/*******************************************************************************
#                        NORTH CAROLINA STATE UNIVERSITY
#
#                              AnyCore Project
# 
# AnyCore written by NCSU authors Rangeen Basu Roy Chowdhury and Eric Rotenberg.
# 
# AnyCore is based on FabScalar which was written by NCSU authors Niket K. 
# Choudhary, Brandon H. Dwiel, and Eric Rotenberg.
# 
# AnyCore also includes contributions by NCSU authors Elliott Forbes, Jayneel 
# Gandhi, Anil Kumar Kannepalli, Sungkwan Ku, Hiran Mayukh, Hashem Hashemi 
# Najaf-abadi, Sandeep Navada, Tanmay Shah, Ashlesha Shastri, Vinesh Srinivasan, 
# and Salil Wadhavkar.
# 
# AnyCore is distributed under the BSD license.
*******************************************************************************/


`timescale 1ns/1ps

//`define PRINT_EN

//`define DUMP_STATS

module simulate();

//* Stop Simulation when COMMIT_COUNT >= SIM_STOP_COUNT
`ifdef SCRATCH_EN
  parameter SIM_STOP_COUNT      = 10_000;
`else
  `ifdef POWER_SIM
    parameter SIM_STOP_COUNT      = 20_000;
  `else
    parameter SIM_STOP_COUNT      = 100_000;
  `endif
`endif

//* Print when (COMMIT_COUNT >= COMMIT_PRINT_COUNT) && (CYCLE_COUNT >= CYCLE_PRINT_COUNT)
parameter COMMIT_PRINT_COUNT  = 0;
parameter CYCLE_PRINT_COUNT   = 0;
parameter STAT_PRINT_COUNT    = 1_000;
parameter IPC_PRINT_COUNT     = 1000;

`ifdef PNR_SIM
  parameter CLKPERIOD           =  100;
`else
  parameter CLKPERIOD           =  `CLKPERIOD;
`endif
parameter IO_CLKPERIOD        =  CLKPERIOD;
//parameter IO_CLKPERIOD        =  CLKPERIOD/20;

`ifdef SCRATCH_EN
  parameter INST_SCRATCH_ENABLED = 1;
  parameter DATA_SCRATCH_ENABLED = 1;
`else
  parameter INST_SCRATCH_ENABLED = 0;
  parameter DATA_SCRATCH_ENABLED = 0;
`endif

`ifdef INST_CACHE
  parameter INST_CACHE_BYPASS = 0;
`else
  parameter INST_CACHE_BYPASS = 1;
`endif

`ifdef DATA_CACHE
  parameter DATA_CACHE_BYPASS = 0;
`else
  parameter DATA_CACHE_BYPASS = 1;
`endif


reg clk_t;
reg clk;
reg ioClk;
reg reset;

reg [5:0] regAddr;
reg [`REG_DATA_WIDTH-1:0] regWrData;
reg [`REG_DATA_WIDTH-1:0] regRdData;
reg       regWrEn;

reg			 data_source; 
reg			 test_mode;   
reg			 data_sourcea;
reg			 test_si1;    
reg			 test_so1;    
reg			 test_si2;    
reg			 test_so2;    
reg			 test_se;    

`ifdef PERF_MON
  reg [`REG_DATA_WIDTH-1:0] perfMonRegAddr; 
  reg [`REG_DATA_WIDTH-1:0] perfMonRegData; 
  reg                       perfMonRegRun ;
  reg                       perfMonRegClr ;
  reg                       perfMonRegGlobalClr ;
`endif

initial
begin
  //$shm_open("waves.shm");
  //$shm_probe(simulate, "ACM");
  //$dumpfile("waves.vcd");
  //$dumpvars(0,fabScalar);
  //$dumplimit(600000000);
end


// Following defines the clk for the simulation.
always #(CLKPERIOD/2.0) 
begin
  clk = ~clk;
end

`ifdef SCAN_EN
  always_comb
  begin
  //  clk =  clk_t & ~test_mode;
    data_source = clk;
  end
`endif
// Following defines the clk for the simulation.
//always #(IO_CLKPERIOD/2.0) 
//begin
//  ioClk = ~ioClk;
//end

always @(*)
  ioClk = clk;

reg  [`SIZE_DATA-1:0]              LOGICAL_REG [`SIZE_RMT-1:0];
reg  [`SIZE_DATA-1:0]              PHYSICAL_REG [`SIZE_PHYSICAL_TABLE-1:0];
reg                                resetFetch;
reg                                verifyCommits;
reg                                cacheModeOverride; //If 1 -> Forces caches to operate in CACHE mode

`ifdef DYNAMIC_CONFIG
  // Power management signals
  reg                                stallFetch;
  reg  [`FETCH_WIDTH-1:0]            fetchLaneActive;
  reg  [`DISPATCH_WIDTH-1:0]         dispatchLaneActive;
  reg  [`ISSUE_WIDTH-1:0]            issueLaneActive;
  reg  [`EXEC_WIDTH-1:0]             execLaneActive;
  reg  [`EXEC_WIDTH-1:0]             saluLaneActive;
  reg  [`EXEC_WIDTH-1:0]             caluLaneActive;
  reg  [`COMMIT_WIDTH-1:0]           commitLaneActive;
  reg  [`NUM_PARTS_RF-1:0]           rfPartitionActive;
  reg  [`NUM_PARTS_RF-1:0]           alPartitionActive;
  reg  [`STRUCT_PARTS_LSQ-1:0]       lsqPartitionActive;
  reg  [`STRUCT_PARTS-1:0]           iqPartitionActive;
  reg  [`STRUCT_PARTS-1:0]           ibuffPartitionActive;
  reg                                reconfigureCore;
`endif

`ifdef SCRATCH_PAD
  reg [`DEBUG_INST_RAM_LOG+`DEBUG_INST_RAM_WIDTH_LOG-1:0]  instScratchAddr;
  reg [7:0]                       instScratchWrData;  
  reg                             instScratchWrEn; 
  reg [`DEBUG_DATA_RAM_LOG+`DEBUG_DATA_RAM_WIDTH_LOG-1:0] dataScratchAddr;
  reg [7:0]                       dataScratchWrData;  
  reg                             dataScratchWrEn;  
  reg [7:0]                       instScratchRdData;  
  reg [7:0]                       dataScratchRdData;  
  reg                             instScratchPadEn = INST_SCRATCH_ENABLED;
  reg                             dataScratchPadEn = DATA_SCRATCH_ENABLED;
`endif

  reg                             instCacheBypass = INST_CACHE_BYPASS;
`ifdef INST_CACHE
  logic [`ICACHE_SIZE_MEM_ADDR-1:0]ic2memReqAddr;     // memory read address
  logic                           ic2memReqValid;     // memory read enable
  logic [`ICACHE_TAG_BITS-1:0]    mem2icTag;          // tag of the incoming data
  logic [`ICACHE_INDEX_BITS-1:0]  mem2icIndex;        // index of the incoming data
  logic [`ICACHE_LINE_SIZE-1:0]   mem2icData;         // requested data
  logic                           mem2icRespValid;    // requested data is ready
`endif  

  logic                              dataCacheBypass = DATA_CACHE_BYPASS;
`ifdef DATA_CACHE
  logic [`DCACHE_SIZE_MEM_ADDR-1:0]  dc2memLdAddr;  // memory read address
  logic                              dc2memLdValid; // memory read enable
  logic [`DCACHE_TAG_BITS-1:0]       mem2dcLdTag;       // tag of the incoming datadetermine
  logic [`DCACHE_INDEX_BITS-1:0]     mem2dcLdIndex;     // index of the incoming data
  logic [`DCACHE_LINE_SIZE-1:0]      mem2dcLdData;      // requested data
  logic                              mem2dcLdValid;     // indicates the requested data is ready
  logic [`DCACHE_SIZE_ST_ADDR-1:0]   dc2memStAddr;  // memory read address
  logic [`SIZE_DATA-1:0]             dc2memStData;  // memory read address
  logic [3:0]                        dc2memStByteEn;  // memory read address
  logic                              dc2memStValid; // memory read enable
  logic                              mem2dcStComplete;
`endif

initial 
begin:INIT_TB
  int i;
//  clk_t                = 0;
  clk                = 0;
  ioClk                = 0;
  reset                = 0;
  regAddr              = 6'h00;
  regWrEn              = 1'b0;
  resetFetch           = 1'b0;
  verifyCommits        = 1'b0;
  cacheModeOverride    = 1'b0;
`ifdef SCAN_EN
  test_mode	       = 1'b1;
`endif
  test_se	       = 1'b0;
`define USE_SDF
  `ifdef USE_SDF
//    `ifdef PNR_SIM
//        $sdf_annotate("../../PNR/out/pr_top_routed.sdf",fab_chip);
//    `else
        $sdf_annotate({"./fab_top.sdf"},fab_chip);
//    `endif
  `endif



  if(!INST_SCRATCH_ENABLED)
  begin
    $initialize_sim();
    $copyMemory();
  end

  $display("");
  $display("");
  $display("**********   ******   ********     *******    ********   ******   ****         ******   ********  ");
  $display("*        *  *      *  *       *   *      *   *       *  *      *  *  *        *      *  *       * ");
  $display("*  ******* *   **   * *  ***   * *   *****  *   ****** *   **   * *  *       *   **   * *  ***   *");
  $display("*  *       *  *  *  * *  *  *  * *  *       *  *       *  *  *  * *  *       *  *  *  * *  *  *  *");
  $display("*  *****   *  ****  * *  ***   * *   ****   *  *       *  ****  * *  *       *  ****  * *  ***   *");
  $display("*      *   *        * *       *   *      *  *  *       *        * *  *       *        * *       * ");
  $display("*  *****   *  ****  * *  ***   *   ****   * *  *       *  ****  * *  *       *  ****  * *  ***   *");
  $display("*  *       *  *  *  * *  *  *  *       *  * *  *       *  *  *  * *  *       *  *  *  * *  *  *  *");
  $display("*  *       *  *  *  * *  ***   *  *****   * *   ****** *  *  *  * *  ******* *  *  *  * *  *  *  *");
  $display("*  *       *  *  *  * *       *   *      *   *       * *  *  *  * *        * *  *  *  * *  *  *  *");
  $display("****       ****  **** ********    *******     ******** ****  **** ********** ****  **** ****  ****");
  $display("");
  $display("FabScalar Copyright (c) 2007-2012 by Niket K. Choudhary, Brandon H. Dwiel, and Eric Rotenberg.");
  $display("All Rights Reserved.");
  $display("");
  $display("");

  if(!INST_SCRATCH_ENABLED)
  begin
    for (i = 0; i < `SIZE_RMT-2; i = i + 1)
    begin
      LOGICAL_REG[i]               = $getArchRegValue(i);
    end

    LOGICAL_REG[32]                = $getArchRegValue(65);
    LOGICAL_REG[33]                = $getArchRegValue(64);

    init_registers();
    $funcsimRunahead();
  end

  clk                            = 0;
  ioClk                          = 0;

`ifdef DYNAMIC_CONFIG  
  stallFetch                     = 1'b0;
  fetchLaneActive                = `FETCH_LANE_ACTIVE     ; 
  dispatchLaneActive             = `DISPATCH_LANE_ACTIVE  ; 
  issueLaneActive                = `ISSUE_LANE_ACTIVE     ; 
  execLaneActive                 = `EXEC_LANE_ACTIVE      ; 
  saluLaneActive                 = `SALU_LANE_ACTIVE      ;
  caluLaneActive                 = `CALU_LANE_ACTIVE      ;
  commitLaneActive               = `COMMIT_LANE_ACTIVE    ; 
  rfPartitionActive              = `RF_PARTITION_ACTIVE   ; 
  alPartitionActive              = `AL_PARTITION_ACTIVE   ; 
  lsqPartitionActive             = `LSQ_PARTITION_ACTIVE  ; 
  iqPartitionActive              = `IQ_PARTITION_ACTIVE   ; 
  ibuffPartitionActive           = `IBUFF_PARTITION_ACTIVE;
  reconfigureCore                = 1'b0;
  
`endif  


  // Assert reset
  #(15*CLKPERIOD) 
  reset                 = 1;
`ifdef SCAN_EN
  stallFetch            = 1'b1;
`endif

  `ifdef PERF_MON
    perfMonRegAddr      = 8'h00;
    perfMonRegClr       = 1'b0;
    perfMonRegRun       = 1'b0;
    perfMonRegGlobalClr = 1'b0;
  `endif

  // Release reset asynchronously to make sure it works
  #(20*CLKPERIOD-4) 
  reset                 = 0;
  #4

  // Let the core run in BIST mode for a while before reconfiguring and loading benchmarks/microkernel
  #(500*CLKPERIOD)

`ifndef SCAN_EN
  stallFetch            = 1'b1;
  #(500*CLKPERIOD)  //Enough time to drain pipeline
  //Reset fetch to start fetching from PC 0x0000 (to load checkpoint and benchmark)
  resetFetch            = 1'b1;
  #(200*CLKPERIOD)  //Enough time to drain pipeline
`endif
  // If in microbenchmark mode, load the kernel and data into scratch pads (or caches)
  if(INST_SCRATCH_ENABLED)
  begin
    // Stall the fetch before loading microbenchmark
  `ifdef DYNAMIC_CONFIG
    #CLKPERIOD
    stallFetch           = 1'b1;  
    #(2*CLKPERIOD)
  `endif

`ifdef SCAN_EN
 //#(2*CLKPERIOD); 
 //data_source = 1'b0;
 #CLKPERIOD; 
 data_sourcea = 1'b0;
 //#(10*CLKPERIOD); 
 //data_source = 1'b1;
 #CLKPERIOD; 
 data_sourcea = 1'b1;
 #(5*CLKPERIOD); 
 data_sourcea = 1'b0;
 scan_in_chain1();
 //scan_out_chain1();
 #(CLKPERIOD) 
 reset                 = 1;
 #(20*CLKPERIOD) 
 reset                 = 0;
 //data_source = 1'b0;
// #50;
 //scan_out_chain1();
 #(20*CLKPERIOD) 
 test_mode = 1'b0;
 //data_source = 1'b0;

//  #(2*CLKPERIOD); 
//  test_mode = 1'b1;
//  data_source = 1'b0;
//  #CLKPERIOD; 
//  data_sourcea = 1'b0;
//  #(10*CLKPERIOD); 
//  data_source = 1'b1;
//  #CLKPERIOD; 
//  data_sourcea = 1'b1;
//  #(5*CLKPERIOD); 
//  data_sourcea = 1'b0;
//  scan_in_chain2();
//  data_source = 1'b0;
 // #50; 
 // scan_out_chain2();
  //test_mode = 1'b0;
`endif
    //$readmemh("kernel.dat",fabScalar.fs1.l1icache.ic.ram);
    //$readmemh("data.dat",fabScalar.lsu.datapath.ldx_path.L1dCache.dc.ram); 
    //for (i = 0; i < 256; i = i + 1)
    //begin
    //    $display("@%d: %08x", i, fabScalar.lsu.datapath.ldx_path.L1dCache.dc.ram[i]);
    //end
 `ifndef SCAN_EN 
    #(200*IO_CLKPERIOD); // Wait for drain to complete
    resetFetch   =   1'b1;
    #(10*IO_CLKPERIOD); // Wait for drain to complete
    load_kernel_scratch();
    read_kernel_scratch();
    load_data_scratch();
    read_data_scratch();
    read_AMT();
    read_PRF();
`endif
    //Unstall the fetch once loading is complete loading microbenchmark
    #(2*CLKPERIOD)
  `ifdef DYNAMIC_CONFIG
    stallFetch           = 1'b0;  
  `endif
  `ifdef SCAN_EN
  #(500*CLKPERIOD)  //Enough time to drain pipeline
  //Reset fetch to start fetching from PC 0x0000 (to load checkpoint and benchmark)
    resetFetch            = 1'b1;
  #(10*CLKPERIOD)
`endif 
    resetFetch           = 1'b0;
    //TODO: Wait for pipeline to be empty
    verifyCommits        = 1'b1;
  end
  // If not in microbenchmark mode, change the cache mode else let it run un SCRATCH mode
  else 
  begin
    stallFetch   =   1'b1;
    #(200*IO_CLKPERIOD); // Wait for drain to complete
    resetFetch   =   1'b1;
    #(10*IO_CLKPERIOD); // Wait for drain to complete
    //load_kernel_scratch();
    //read_kernel_scratch();
    //load_data_scratch();
    //read_data_scratch();
    //read_AMT();
    //read_PRF();
 
    // Test the cache mode override
    cacheModeOverride = 1'b1;

    #(5*CLKPERIOD)
    //TODO: Wait for pipeline to be empty
    verifyCommits        = 1'b1;
    stallFetch           = 1'b0;
    resetFetch           = 1'b0;
    #(2*CLKPERIOD)
    // If not in microbenchmark mode, let the core run in CACHE mode for a while with actual 
    // benchmark before reconfiguring
    #(1000*CLKPERIOD)
    verifyCommits        = 1'b1; // Dummy statement to avoid error. Doesn't really do anything
  end


//load_checkpoint_PRF();
//read_checkpoint_PRF();
  
`ifdef DYNAMIC_CONFIG


  // Stall the fetch before reconfiguring
  // TODO: Test that it works without this as well
  #CLKPERIOD
`ifdef SCAN_EN
  #(10000*CLKPERIOD)
`endif 
  stallFetch           = 1'b1;  

  #(10*IO_CLKPERIOD)

  regWrEn     = 1'b0;
  regAddr     = 6'h01;
  regWrData   = {{(`REG_DATA_WIDTH-`FETCH_WIDTH){1'b0}},fetchLaneActive}     ; 
  regWrEn     = 1'b1;
  #IO_CLKPERIOD
  regWrEn     = 1'b0;
  #IO_CLKPERIOD
  regAddr     = 6'h02;
  regWrData   = {{(`REG_DATA_WIDTH-`DISPATCH_WIDTH){1'b0}},dispatchLaneActive}     ; 
  regWrEn     = 1'b1;
  #IO_CLKPERIOD
  regWrEn     = 1'b0;
  #IO_CLKPERIOD
  regAddr     = 6'h03;
  regWrData   = {{(`REG_DATA_WIDTH-`ISSUE_WIDTH){1'b0}},issueLaneActive}     ; 
  regWrEn     = 1'b1;
  #IO_CLKPERIOD
  regWrEn     = 1'b0;
  #IO_CLKPERIOD
  regAddr     = 6'h04;
  regWrData   = {{(`REG_DATA_WIDTH-`EXEC_WIDTH){1'b0}},execLaneActive}     ; 
  regWrEn     = 1'b1;
  #IO_CLKPERIOD
  regWrEn     = 1'b0;
  #IO_CLKPERIOD
  regAddr     = 6'h05;
  regWrData   = {{(`REG_DATA_WIDTH-`EXEC_WIDTH){1'b0}},saluLaneActive}     ; 
  regWrEn     = 1'b1;
  #IO_CLKPERIOD
  regWrEn     = 1'b0;
  #IO_CLKPERIOD
  regAddr     = 6'h06;
  regWrData   = {{(`REG_DATA_WIDTH-`EXEC_WIDTH){1'b0}},caluLaneActive}     ; 
  regWrEn     = 1'b1;
  #IO_CLKPERIOD
  regWrEn     = 1'b0;
  #IO_CLKPERIOD
  regAddr     = 6'h07;
  regWrData   = {{(`REG_DATA_WIDTH-`COMMIT_WIDTH){1'b0}},commitLaneActive}     ; 
  regWrEn     = 1'b1;
  #IO_CLKPERIOD
  regWrEn     = 1'b0;
  #IO_CLKPERIOD
  regAddr     = 6'h08;
  regWrData   = {{`REG_DATA_WIDTH-`NUM_PARTS_RF{1'b0}},rfPartitionActive}     ; 
  regWrEn     = 1'b1;
  #IO_CLKPERIOD
  regWrEn     = 1'b0;
  #IO_CLKPERIOD
  regAddr     = 6'h09;
  regWrData   = {{`REG_DATA_WIDTH-`NUM_PARTS_RF{1'b0}},alPartitionActive}     ; 
  regWrEn     = 1'b1;
  #IO_CLKPERIOD
  regWrEn     = 1'b0;
  #IO_CLKPERIOD
  regAddr     = 6'h0A;
  regWrData   = {{`REG_DATA_WIDTH-`STRUCT_PARTS{1'b0}},lsqPartitionActive}     ; 
  regWrEn     = 1'b1;
  #IO_CLKPERIOD
  regWrEn     = 1'b0;
  #IO_CLKPERIOD
  regAddr     = 6'h0B;
  regWrData   = {{`REG_DATA_WIDTH-`STRUCT_PARTS{1'b0}},iqPartitionActive}     ; 
  regWrEn     = 1'b1;
  #IO_CLKPERIOD
  regWrEn     = 1'b0;
  #IO_CLKPERIOD
  regAddr     = 6'h0C;
  regWrData   = {{`REG_DATA_WIDTH-`STRUCT_PARTS{1'b0}},ibuffPartitionActive}     ; 
  regWrEn     = 1'b1;
  #IO_CLKPERIOD
  regWrEn     = 1'b0;
  #IO_CLKPERIOD


  /* Post reconfiguration reset sequence*/
  #(IO_CLKPERIOD)
  reconfigureCore      = 1'b1;
  #(20*IO_CLKPERIOD)
  reconfigureCore      = 1'b0;

  // Unstall the fetch
  #IO_CLKPERIOD
  stallFetch           = 1'b0;
  #(1000*IO_CLKPERIOD)

  //Change mode of the caches to CACHE mode
  regWrEn     = 1'b0;
  regAddr     = 6'h1F;
  regWrData   = 8'b00000000     ; //00 is cache mode 
  regWrEn     = 1'b1;
  #IO_CLKPERIOD
  regWrEn     = 1'b0;


`ifdef SCRATCH_EN  
  // Disable the scratch pads
  regAddr     = 6'h0D; 
  regWrData   = 8'h0;
  regWrEn     = 1'b1;
  #IO_CLKPERIOD
  regWrEn     = 1'b0;
`endif

  // Deassert the override and let the normal
  // config take effect.
  #(100*IO_CLKPERIOD)
  cacheModeOverride = 1'b0;

`endif 

end


reg  [`SIZE_PC-1:0]                instPC_tb [0:`FETCH_WIDTH-1];
reg  [`SIZE_PC-1:0]                instPC;
wire [`ICACHE_PC_PKT_BITS-1:0]     instPC_packet;
wire [`ICACHE_INST_PKT_BITS-1:0]   inst_packet;
reg  [`SIZE_INSTRUCTION-1:0]       inst_tb   [0:`FETCH_WIDTH-1];
reg  [`FETCH_WIDTH*`SIZE_INSTRUCTION-1:0]       inst;

wire [`SIZE_PC-1:0]                memAddr;

wire [`SIZE_PC-1:0]                ldAddr;
wire [`SIZE_DATA-1:0]              ldData;
wire                               ldEn;

wire [`SIZE_PC-1:0]                stAddr;
wire [`SIZE_DATA-1:0]              stData;
wire [3:0]                         stEn;

reg [`SIZE_DATA_BYTE_OFFSET+`SIZE_PHYSICAL_LOG-1:0] debugPRFAddr  ;
reg [`SRAM_DATA_WIDTH-1:0] 			   debugPRFWrData;             
reg 					                     debugPRFWrEn  = 1'b0;
reg [`SRAM_DATA_WIDTH-1:0] 			   debugPRFRdData;

wire [`SIZE_PC-1:0]                ldAddr_tmp;
wire [`DCACHE_LD_ADDR_PKT_BITS-1:0]ldAddr_packet;
wire [`DCACHE_LD_DATA_PKT_BITS-1:0]ldData_packet;

wire [`SIZE_PC-1:0]                stAddr_tmp;
wire [`SIZE_DATA-1:0]              stData_tmp;
wire [3:0]                         stEn_tmp;
wire [`DCACHE_ST_PKT_BITS-1:0]     st_packet;


`ifdef PNR_SIM
  pr_top fab_chip();
  
assign fab_chip.pi_any_regAddr_i_0.P        = regAddr[0]; 
assign fab_chip.pi_any_regAddr_i_1.P        = regAddr[1]; 
assign fab_chip.pi_any_regAddr_i_2.P        = regAddr[2]; 
assign fab_chip.pi_any_regAddr_i_3.P        = regAddr[3]; 
assign fab_chip.pi_any_regAddr_i_4.P        = regAddr[4]; 
assign fab_chip.pi_any_regAddr_i_5.P        = regAddr[5]; 
assign fab_chip.pi_any_regWrData_i_0.P      = regWrData[0]; 
assign fab_chip.pi_any_regWrData_i_1.P      = regWrData[1]; 
assign fab_chip.pi_any_regWrData_i_2.P      = regWrData[2]; 
assign fab_chip.pi_any_regWrData_i_3.P      = regWrData[3]; 
assign fab_chip.pi_any_regWrData_i_4.P      = regWrData[4]; 
assign fab_chip.pi_any_regWrData_i_5.P      = regWrData[5]; 
assign fab_chip.pi_any_regWrData_i_6.P      = regWrData[6]; 
assign fab_chip.pi_any_regWrData_i_7.P      = regWrData[7]; 
assign fab_chip.pi_any_reconfigureCore_i.P  = reconfigureCore; 
assign fab_chip.pi_any_inst_packet_i_0.P    = inst_packet[0]; 
assign fab_chip.pi_any_inst_packet_i_1.P    = inst_packet[1]; 
assign fab_chip.pi_any_inst_packet_i_2.P    = inst_packet[2]; 
assign fab_chip.pi_any_inst_packet_i_3.P    = inst_packet[3]; 
assign fab_chip.pi_any_inst_packet_i_4.P    = inst_packet[4]; 
assign fab_chip.pi_any_inst_packet_i_5.P    = inst_packet[5]; 
assign fab_chip.pi_any_inst_packet_i_6.P    = inst_packet[6]; 
assign fab_chip.pi_any_inst_packet_i_7.P    = inst_packet[7]; 
assign fab_chip.pi_any_clk.P                = clk; 
assign fab_chip.pi_any_reset.P              = reset;
assign fab_chip.pi_any_mem2dcStComplete_i.P = mem2dcStComplete;
assign fab_chip.pi_any_ldData_packet_i_0.P  = ldData_packet[0]; 
assign fab_chip.pi_any_ldData_packet_i_1.P  = ldData_packet[1]; 
assign fab_chip.pi_any_ldData_packet_i_2.P  = ldData_packet[2]; 
assign fab_chip.pi_any_ldData_packet_i_3.P  = ldData_packet[3]; 
assign fab_chip.pi_any_ldData_packet_i_4.P  = ldData_packet[4]; 
assign fab_chip.pi_any_ldData_packet_i_5.P  = ldData_packet[5]; 
assign fab_chip.pi_any_ldData_packet_i_6.P  = ldData_packet[6]; 
assign fab_chip.pi_any_ldData_packet_i_7.P  = ldData_packet[7]; 
assign fab_chip.pi_any_regWrEn_i.P          = regWrEn; 
assign fab_chip.pi_any_stallFetch_i.P       = stallFetch;
assign fab_chip.pi_any_data_source.P        = 1'b0;
assign fab_chip.pi_any_test_mode.P          = 1'b0;
assign fab_chip.pi_any_data_sourcea.P       = 1'b0;
assign fab_chip.pi_any_test_si1.P           = 1'bx;
assign fab_chip.pi_any_test_si2.P           = 1'bx;
assign fab_chip.pi_any_test_se.P            = 1'b0;
assign fab_chip.pi_any_resetFetch_i.P       = resetFetch; 
assign fab_chip.pi_any_cacheModeOverride_i.P= cacheModeOverride;


//assign  = fab_chip/po_any_test_so1.P      ; 
//assign  = fab_chip/po_any_test_so2.P      ; 
assign  regRdData[0]      = fab_chip.po_any_regRdData_o_0.P      ; 
assign  regRdData[1]      = fab_chip.po_any_regRdData_o_1.P      ; 
assign  regRdData[2]      = fab_chip.po_any_regRdData_o_2.P      ; 
assign  regRdData[3]      = fab_chip.po_any_regRdData_o_3.P      ; 
assign  regRdData[4]      = fab_chip.po_any_regRdData_o_4.P      ; 
assign  regRdData[5]      = fab_chip.po_any_regRdData_o_5.P      ; 
assign  regRdData[6]      = fab_chip.po_any_regRdData_o_6.P      ; 
assign  regRdData[7]      = fab_chip.po_any_regRdData_o_7.P      ; 
assign  instPC_packet[0]  = fab_chip.po_any_instPC_packet_o_0.P      ; 
assign  instPC_packet[1]  = fab_chip.po_any_instPC_packet_o_1.P      ; 
assign  instPC_packet[2]  = fab_chip.po_any_instPC_packet_o_2.P      ; 
assign  instPC_packet[3]  = fab_chip.po_any_instPC_packet_o_3.P      ; 
assign  instPC_packet[4]  = fab_chip.po_any_instPC_packet_o_4.P      ; 
assign  instPC_packet[5]  = fab_chip.po_any_instPC_packet_o_5.P      ; 
assign  instPC_packet[6]  = fab_chip.po_any_instPC_packet_o_6.P      ; 
assign  instPC_packet[7]  = fab_chip.po_any_instPC_packet_o_7.P      ; 
assign  st_packet[0]      = fab_chip.po_any_st_packet_o_0.P      ; 
assign  st_packet[1]      = fab_chip.po_any_st_packet_o_1.P      ; 
assign  st_packet[2]      = fab_chip.po_any_st_packet_o_2.P      ; 
assign  st_packet[3]      = fab_chip.po_any_st_packet_o_3.P      ; 
assign  st_packet[4]      = fab_chip.po_any_st_packet_o_4.P      ; 
assign  st_packet[5]      = fab_chip.po_any_st_packet_o_5.P      ; 
assign  st_packet[6]      = fab_chip.po_any_st_packet_o_6.P      ; 
assign  st_packet[7]      = fab_chip.po_any_st_packet_o_7.P      ; 
assign  ldAddr_packet[0]  = fab_chip.po_any_ldAddr_packet_o_0.P      ; 
assign  ldAddr_packet[1]  = fab_chip.po_any_ldAddr_packet_o_1.P      ; 
assign  ldAddr_packet[2]  = fab_chip.po_any_ldAddr_packet_o_2.P      ; 
assign  ldAddr_packet[3]  = fab_chip.po_any_ldAddr_packet_o_3.P      ; 
assign  ldAddr_packet[4]  = fab_chip.po_any_ldAddr_packet_o_4.P      ; 
assign  ldAddr_packet[5]  = fab_chip.po_any_ldAddr_packet_o_5.P      ; 
assign  ldAddr_packet[6]  = fab_chip.po_any_ldAddr_packet_o_6.P      ; 
assign  ldAddr_packet[7]  = fab_chip.po_any_ldAddr_packet_o_7.P      ; 
assign  toggleFlag        = fab_chip.po_any_toggleFlag_o.P      ; 

`else
  fab_top fab_chip(
  
      .clk                                 (clk),
      //.coreClk                             (clk),
      //.ioClk                               (ioClk),
      .reset                               (reset),
      .resetFetch_i                        (resetFetch),
      .cacheModeOverride_i                 (cacheModeOverride),
      .toggleFlag_o                        (toggleFlag),

 `ifndef SCAN_EN 
      .data_source                         (1'b0), 
      .test_mode                           (1'b0),
      .data_sourcea                        (1'b0), 
      .test_si1                            (), 
      .test_so1                            (), 
      .test_si2                            (), 
      .test_so2                            (), 
      .test_se                             (1'b0),
`else
     .data_source                         (data_source), 
     .test_mode                           (test_mode),
     .data_sourcea                        (data_sourcea), 
     .test_si1                            (test_si1), 
     .test_so1                            (test_so1), 
     .test_si2                            (test_si2), 
     .test_so2                            (test_so2), 
     .test_se                             (test_se),
`endif 
      .regAddr_i                           (regAddr),
      .regWrData_i                         (regWrData),
      .regWrEn_i                           (regWrEn),
      .regRdData_o                         (regRdData),
  
      .stallFetch_i                        (stallFetch),
      .reconfigureCore_i                   (reconfigureCore),
  
      /* Parallel interface for debug and simulation only */
      /* To instruction memory */
      //.instPC_o                            (instPC),
      //.inst_i                              (inst),
  
  	  /* To data memory */
      //.ldAddr_o                            (ldAddr),
      //.ldData_i                            (ldData),
      //.ldEn_o                              (ldEn),
  
      //.stAddr_o                            (stAddr),
      //.stData_o                            (stData),
      //.stEn_o                              (stEn),
      /* Parallel interface ends */
  
    `ifdef DATA_CACHE
      .mem2dcStComplete_i                 (mem2dcStComplete),
    `endif
  
  
      /* Packet interface for fabrication */
      // Operates at ioClk
      .instPC_packet_o                     (instPC_packet),
      .inst_packet_i                       (inst_packet),
  
      .ldAddr_packet_o                     (ldAddr_packet),
      .ldData_packet_i                     (ldData_packet),
      .st_packet_o                         (st_packet)
      /* Packet interface ends */
  
   );
`endif

`ifdef INST_CACHE

  logic [32-`ICACHE_SIZE_MEM_ADDR-1:0] instDePktDummy;
  
  Depacketizer #(
      .PAYLOAD_WIDTH      (32),
      .PACKET_WIDTH       (`ICACHE_PC_PKT_BITS),
      .ID                 (0),
      .DEPTH              (4),
      .DEPTH_LOG          (2),
      .N_PKTS_BITS        (2),
      .INST_NAME          ("instPC_depkt_tb")
  )
      instPC_depacketizer (
  
      .reset              (reset),
  
      .clk_packet         (ioClk),
      .packet_i           (instPC_packet),
      .packet_af_o        (instPC_depacket_af),
  
      .clk_payload        (ioClk),
      .payload_o          ({instDePktDummy,ic2memReqAddr}),
      .payload_valid_o    (ic2memReqValid),
      .packet_received_o  ()
  );
  
  logic [32-`ICACHE_SIZE_MEM_ADDR-1:0] instPktDummy = {(32-`ICACHE_SIZE_MEM_ADDR){1'b0}};
  
  Packetizer_wide #(
      .PAYLOAD_WIDTH          (32+`ICACHE_LINE_SIZE),
      .PACKET_WIDTH           (`ICACHE_INST_PKT_BITS),
      .ID                     (1),
      .DEPTH                  (4),
      .DEPTH_LOG              (2),
      .N_PKTS_BITS            (2),
      .THROTTLE               (0) //Throttling is disabled
  )
      inst_packetizer (
  
      .reset                  (reset),
  
      .clk_payload            (ioClk),
      .payload_req_i          (mem2icRespValid), //Looped back from Depacketizer
      .payload_i              ({instPktDummy,mem2icTag,mem2icIndex,mem2icData}),
      .payload_grant_o        (),
      .push_af_o              (inst_push_af),
  
      .clk_packet             (ioClk),
      .packet_req_o           (inst_packet_req),
      .lock_o                 (),
      .packet_o               (inst_packet),
      .packet_grant_i         (inst_packet_req), //Request is looped back in as grant
      .packet_received_i      (1'b0)
  );
`endif //ifdef INST_CACHE

`ifdef DATA_CACHE

  logic [32-`DCACHE_SIZE_MEM_ADDR-1:0] ldDePktDummy;

  Depacketizer #(
      .PAYLOAD_WIDTH      (32),
      .PACKET_WIDTH       (`DCACHE_LD_ADDR_PKT_BITS),
      .ID                 (0),
      .DEPTH              (4),
      .DEPTH_LOG          (2),
      .N_PKTS_BITS        (2),
      .INST_NAME          ("ldAddr_depkt_tb")
  )
      ldAddr_depacketizer (
  
      .reset              (reset),
  
      .clk_packet         (ioClk),
      .packet_i           (ldAddr_packet),
      .packet_af_o        (ldAddr_depacket_af),
  
      .clk_payload        (ioClk),
      //.payload_o          (ldAddr_tmp),
      .payload_o          ({ldDePktDummy,dc2memLdAddr}),
      .payload_valid_o    (dc2memLdValid),
      .packet_received_o  ()
  );
  
  logic [32-`DCACHE_SIZE_MEM_ADDR-1:0] ldPktDummy = {(32-`DCACHE_SIZE_MEM_ADDR){1'b0}};
  
  Packetizer #(
      .PAYLOAD_WIDTH          (32+`DCACHE_LINE_SIZE),
      .PACKET_WIDTH           (`DCACHE_LD_DATA_PKT_BITS),
      .ID                     (1),
      .DEPTH                  (4),
      .DEPTH_LOG              (2),
      .N_PKTS_BITS            (2),
      .THROTTLE               (0) //Throttling is disabled
  )
      ldData_packetizer (
  
      .reset                  (reset),
  
      .clk_payload            (ioClk),
      .payload_req_i          (mem2dcLdValid),
      .payload_i              ({ldPktDummy,mem2dcLdTag,mem2dcLdIndex,mem2dcLdData}),
      .payload_grant_o        (),
      .push_af_o              (ldData_push_af),
  
      .clk_packet             (ioClk),
      .packet_req_o           (ldData_packet_req),
      .lock_o                 (),
      .packet_o               (ldData_packet),
      .packet_grant_i         (ldData_packet_req), //Request is looped back in as grant
      .packet_received_i      (1'b0)
  );
  
  
  
  logic [36-`DCACHE_SIZE_ST_ADDR-1:0] stDePktDummy;
  
  Depacketizer #(
      .PAYLOAD_WIDTH      (4+32+32+4),
      .PACKET_WIDTH       (`DCACHE_ST_PKT_BITS),
      .ID                 (0),
      .DEPTH              (4),
      .DEPTH_LOG          (2),
      .N_PKTS_BITS        (2),
      .INST_NAME          ("st_depkt_tb")
  )
      st_depacketizer (
  
      .reset              (reset),
  
      .clk_packet         (ioClk),
      .packet_i           (st_packet),
      .packet_af_o        (st_depacket_af),
  
      .clk_payload        (ioClk),
      .payload_o          ({stDePktDummy,dc2memStAddr,dc2memStData,dc2memStByteEn}),
      .payload_valid_o    (dc2memStValid),
      .packet_received_o  ()
  );
`endif //ifdef DATA_CACHE


//assign  ldAddr = memAddr;
//assign  stAddr = memAddr;
always_comb
begin:INST_PC
  int i;
  for(i = 0;i < `FETCH_WIDTH; i++)
  begin
    instPC_tb[i] = instPC+(8*i);
    inst[((i+1)*`SIZE_INSTRUCTION-1)-:`SIZE_INSTRUCTION] = inst_tb[i];
  end
end

memory_hier mem (
    .icClk                               (ioClk),
    .dcClk                               (ioClk),
    .reset                               (reset),

    .icPC_i                              (instPC_tb),
    .icInstReq_i                         (instReq & (INST_SCRATCH_ENABLED ? 1'b0 : 1'b1)), //Mask requests to prevent crash
    .icInst_o                            (inst_tb),

  `ifdef INST_CACHE
    .ic2memReqAddr_i                     (ic2memReqAddr),
    .ic2memReqValid_i                    (ic2memReqValid & (INST_SCRATCH_ENABLED ? 1'b0 : 1'b1)), //Mask requests to prevent crash
    .mem2icTag_o                         (mem2icTag), 
    .mem2icIndex_o                       (mem2icIndex),     
    .mem2icData_o                        (mem2icData),      
    .mem2icRespValid_o                   (mem2icRespValid), 
  `endif

  `ifdef DATA_CACHE
    .dc2memLdAddr_i                      (dc2memLdAddr     ), // memory read address
    .dc2memLdValid_i                     (dc2memLdValid  & (DATA_SCRATCH_ENABLED ? 1'b0 : 1'b1)), // memory read enable
                                                            
    .mem2dcLdTag_o                       (mem2dcLdTag      ), // tag of the incoming datadetermine
    .mem2dcLdIndex_o                     (mem2dcLdIndex    ), // index of the incoming data
    .mem2dcLdData_o                      (mem2dcLdData     ), // requested data
    .mem2dcLdValid_o                     (mem2dcLdValid    ), // indicates the requested data is ready
                                                            
    .dc2memStAddr_i                      (dc2memStAddr     ), // memory read address
    .dc2memStData_i                      (dc2memStData     ), // memory read address
    .dc2memStByteEn_i                    (dc2memStByteEn   ), // memory read address
    .dc2memStValid_i                     (dc2memStValid  & (DATA_SCRATCH_ENABLED ? 1'b0 : 1'b1)), // memory read enable
                                                            
    .mem2dcStComplete_o                  (mem2dcStComplete ),
  `endif    
  
    .ldAddr_i                            (ldAddr),
    .ldData_o                            (ldData),
    .ldEn_i                              (ldEn  & (DATA_SCRATCH_ENABLED ? 1'b0 : 1'b1)),

    .stAddr_i                            (stAddr),
    .stData_i                            (stData),
    .stEn_i                              (stEn & (DATA_SCRATCH_ENABLED ? 4'b0000 : 4'b1111))
);

integer CYCLE_COUNT;
integer COMMIT_COUNT;

/*
always @(posedge clk)
begin:HANDLE_EXCEPTION
  int i;
  reg [`SIZE_PC-1:0] TRAP_PC;
  if(!INST_SCRATCH_ENABLED) // This is controlled in the testbench
  begin

  // Following code handles the SYSCALL (trap).
  if (fab_chip.fabScalar.activeList.exceptionFlag[0] && (|fab_chip.fabScalar.activeList.alCount))
  begin

    //Functional simulator is stalled waiting to execute the trap.
    //Signal it to proceed with the trap.
    

    TRAP_PC = fab_chip.fabScalar.activeList.commitPC[0];

      $display("TRAP (Cycle: %0d PC: %08x Code: %0d)\n",
               CYCLE_COUNT,
               TRAP_PC,
               $getArchRegValue(2));

      if ($getArchRegValue(2) == 1)
      begin
          $display("SS_SYS_exit encountered. Exiting the simulation");
          $finish;
      end

      $handleTrap();

      //The memory state of the timing simulator is now stale.
      //Copy values from the functional simulator.
      
      $copyMemory();

      //Registers of the timing simulator are now stale.
      //Copy values from the functional simulator.
      
      for (i = 0; i < `SIZE_RMT - 2; i++) 
      begin
        LOGICAL_REG[i]  = $getArchRegValue(i);
      end

      LOGICAL_REG[32]   = $getArchRegValue(65);
      LOGICAL_REG[33]   = $getArchRegValue(64);

      //Functional simulator is waiting to resume after the trap.
      //Signal it to resume.
      
      $resumeTrap();

      $getRetireInstPC(1,CYCLE_COUNT,TRAP_PC,0,0,0);
      init_registers;
    end
  end // !INST_SCRATCH_ENABLED

  //After the SYSCALL is handled by the functional simulator, architectural
  //values from functional simulator should be copied to the Register File.
  
  if (fab_chip.fabScalar.activeList.exceptionFlag_reg) 
  begin
    $display("CYCLE:%d Exception is High\n", CYCLE_COUNT);
    // init_registers; 
    // copyRF; 
    // copySimRF; 
  end
end
*/

reg [3:0]                    totalCommit;
wire    PRINT;
assign  PRINT = (COMMIT_COUNT >= COMMIT_PRINT_COUNT) && (CYCLE_COUNT > CYCLE_PRINT_COUNT);

integer last_commit_cnt;
integer load_violation_count;
integer br_count;
integer br_mispredict_count;
integer ld_count;
integer btb_miss;
integer btb_miss_rtn;
integer fetch1_stall;
integer ctiq_stall;
integer instBuf_stall;
integer freelist_stall;
integer smt_stall;
integer backend_stall;
integer rob_stall;
integer iq_stall;
integer ldq_stall;
integer stq_stall;

// cti stats ////////////////////
`define     stat_num_corr           fab_chip.fabScalar.exePipe1.execute.stat_num_corr
`define     stat_num_pred           fab_chip.fabScalar.exePipe1.execute.stat_num_pred
`define     stat_num_cond_corr      fab_chip.fabScalar.exePipe1.execute.stat_num_cond_corr
`define     stat_num_cond_pred      fab_chip.fabScalar.exePipe1.execute.stat_num_cond_pred
`define     stat_num_return_corr    fab_chip.fabScalar.exePipe1.execute.stat_num_return_corr
`define     stat_num_return_pred    fab_chip.fabScalar.exePipe1.execute.stat_num_return_pred
/////////////////////////////////

int     ib_count;
int     fl_count;
int     iq_count;
int     ldq_count;
int     stq_count;
int     al_count;

int     commit_1;
int     commit_2;
int     commit_3;
int     commit_4;

real    ib_avg;
real    fl_avg;
real    iq_avg;
real    ldq_avg;
real    stq_avg;
real    al_avg;

real    ipc;

integer fd0;
integer fd1;
integer fd2;
integer fd3;
integer fd4;
integer fd5;
integer fd6;
integer fd7;
integer fd8;
integer fd9;
integer fd10;
integer fd11;
integer fd12;
integer fd13;
integer fd14;
integer fd16;
integer fd17;
integer fd18;
integer fd19;
integer fd20;
integer fd21;
integer fd22;
integer fd23;

initial
begin
    CYCLE_COUNT          = 0;
    COMMIT_COUNT         = 0;
    load_violation_count = 0;
    br_count             = 0;
    br_mispredict_count  = 0;
    ld_count             = 0;
    btb_miss             = 0;
    btb_miss_rtn         = 0;
    fetch1_stall         = 0;
    ctiq_stall           = 0;
    instBuf_stall        = 0;
    freelist_stall       = 0;
    smt_stall            = 0;
    backend_stall        = 0;
    rob_stall            = 0;
    iq_stall             = 0;
    ldq_stall            = 0;
    stq_stall            = 0;
    last_commit_cnt      = 0;

    ib_count             = 0;
    fl_count             = 0;
    iq_count             = 0;
    ldq_count            = 0;
    stq_count            = 0;
    al_count             = 0;

    commit_1             = 0;
    commit_2             = 0;
    commit_3             = 0;
    commit_4             = 0;

    fd9         = $fopen("results/fetch1.txt","w");
    fd14        = $fopen("results/fetch2.txt","w");
    fd2         = $fopen("results/decode.txt","w");
    fd1         = $fopen("results/instBuf.txt","w");
    fd0         = $fopen("results/rename.txt","w");
    fd3         = $fopen("results/dispatch.txt","w");
    fd4         = $fopen("results/select.txt","w");
    fd5         = $fopen("results/issueq.txt","w");
    fd6         = $fopen("results/regread.txt","w");
    fd23        = $fopen("results/PhyRegFile.txt","w");
    fd13        = $fopen("results/exe.txt","w");
    fd7         = $fopen("results/activeList.txt","w");
    fd10        = $fopen("results/lsu.txt","w");
    fd8         = $fopen("results/writebk.txt","w");

    fd16        = $fopen("results/statistics.txt","w");
    fd17        = $fopen("results/fabscalar.txt","w");

`ifdef DUMP_STATS
    $fwrite(fd16, "CYCLE, "); 
    $fwrite(fd16, "COMMIT, "); 

    $fwrite(fd16, "IB-avg, "); 
    $fwrite(fd16, "FL-avg, "); 
    $fwrite(fd16, "IQ-avg, "); 
    $fwrite(fd16, "LDQ-avg, "); 
    $fwrite(fd16, "STQ-avg, "); 
    $fwrite(fd16, "AL-avg, "); 

    $fwrite(fd16, "FS1-stall, ");
    $fwrite(fd16, "CTI-stall, ");
    $fwrite(fd16, "IB-stall, ");
    $fwrite(fd16, "FL-stall, ");
    $fwrite(fd16, "BE-stall, ");
    $fwrite(fd16, "LDQ-stall, ");
    $fwrite(fd16, "STQ-stall, ");
    $fwrite(fd16, "IQ-stall, ");
    $fwrite(fd16, "AL-stall, ");

    $fwrite(fd16, "BTB-Miss, ");
    $fwrite(fd16, "Miss-Rtn, ");
    $fwrite(fd16, "BR-Count, ");
    $fwrite(fd16, "Mis-Cnt, ");
    $fwrite(fd16, "LdVio-Cnt, ");

    $fwrite(fd16, "stat_num_corr, ");
    $fwrite(fd16, "stat_num_pred, ");
    $fwrite(fd16, "stat_num_cond_corr, ");
    $fwrite(fd16, "stat_num_cond_pred, ");
    $fwrite(fd16, "stat_num_return_corr, ");
    $fwrite(fd16, "stat_num_return_pred, ");

    $fwrite(fd16, "Commit_1, ");
    $fwrite(fd16, "Commit_2, ");
    $fwrite(fd16, "Commit_3, ");
    $fwrite(fd16, "Commit_4\n");
`endif
end


always @(posedge clk)
begin: HEARTBEAT
    
    CYCLE_COUNT = CYCLE_COUNT + 1;

    COMMIT_COUNT = COMMIT_COUNT + totalCommit;

    if ((CYCLE_COUNT % STAT_PRINT_COUNT) == 0)
    begin
        if (((COMMIT_COUNT - last_commit_cnt) == 0) & verifyCommits) // Check for stalls only once benchmark has started
        begin
            $display("Cycle Count:%d Commit Count:%d  BTB-Miss:%d BTB-Miss-Rtn:%d  Br-Count:%d Br-Mispredict:%d",
                     CYCLE_COUNT,
                     COMMIT_COUNT,
                     btb_miss,
                     btb_miss_rtn,
                     br_count,
                     br_mispredict_count);

            $display("ERROR: instruction committing has stalled (Cycle: %0d, Commit: %0d", CYCLE_COUNT, COMMIT_COUNT);
            $finish;
            read_AMT();
            read_PRF();
          `ifdef PERF_MON
            read_perf_mon();
          `endif  


        end

        $display("Cycle: %d Commit: %d  BTB-Miss: %0d  BTB-Miss-Rtn: %0d  Br-Count: %0d  Br-Mispredict: %0d",
                 CYCLE_COUNT,
                 COMMIT_COUNT,
                 btb_miss,
                 btb_miss_rtn,
                 br_count,
                 br_mispredict_count);

        
`ifdef DUMP_STATS
        ib_avg    = ib_count/(CYCLE_COUNT-10.0);
        fl_avg    = fl_count/(CYCLE_COUNT-10.0);
        iq_avg    = iq_count/(CYCLE_COUNT-10.0);
        ldq_avg   = ldq_count/(CYCLE_COUNT-10.0);
        stq_avg   = stq_count/(CYCLE_COUNT-10.0);
        al_avg    = al_count/(CYCLE_COUNT-10.0);

        $fwrite(fd16, "%d, ", CYCLE_COUNT); 
        $fwrite(fd16, "%d, ", COMMIT_COUNT); 

        $fwrite(fd16, "%2.3f, ", ib_avg); 
        $fwrite(fd16, "%2.3f, ", fl_avg); 
        $fwrite(fd16, "%2.3f, ", iq_avg); 
        $fwrite(fd16, "%2.4f, ", ldq_avg); 
        $fwrite(fd16, "%2.4f, ", stq_avg); 
        $fwrite(fd16, "%2.3f, ", al_avg); 

        $fwrite(fd16, "%d, ", fetch1_stall); 
        $fwrite(fd16, "%d, ", ctiq_stall); 
        $fwrite(fd16, "%d, ", instBuf_stall); 
        $fwrite(fd16, "%d, ", freelist_stall); 
        $fwrite(fd16, "%d, ", backend_stall); 
        $fwrite(fd16, "%d, ", ldq_stall); 
        $fwrite(fd16, "%d, ", stq_stall); 
        $fwrite(fd16, "%d, ", iq_stall); 
        $fwrite(fd16, "%d, ", rob_stall); 

        $fwrite(fd16, "%d, ", btb_miss); 
        $fwrite(fd16, "%d, ", btb_miss_rtn); 
        $fwrite(fd16, "%d, ", br_count); 
        $fwrite(fd16, "%d, ", br_mispredict_count); 
        $fwrite(fd16, "%d, ", load_violation_count); 

        $fwrite(fd16, "%d, ", `stat_num_corr);
        $fwrite(fd16, "%d, ", `stat_num_pred);
        $fwrite(fd16, "%d, ", `stat_num_cond_corr);
        $fwrite(fd16, "%d, ", `stat_num_cond_pred);
        $fwrite(fd16, "%d, ", `stat_num_return_corr);
        $fwrite(fd16, "%d, ", `stat_num_return_pred);

        $fwrite(fd16, "%d, ", commit_1); 
        $fwrite(fd16, "%d, ", commit_2); 
        $fwrite(fd16, "%d, ", commit_3); 
        $fwrite(fd16, "%d\n", commit_4); 
`endif

        last_commit_cnt = COMMIT_COUNT;
    end
end
/*
fuPkt                           exePacket      [0:`ISSUE_WIDTH-1];

always_comb
begin

    exePacket[0]      = fab_chip.fabScalar.exePipe0.exePacket;
    exePacket[1]      = fab_chip.fabScalar.exePipe1.exePacket;
    exePacket[2]      = fab_chip.fabScalar.exePipe2.exePacket;
`ifdef ISSUE_FOUR_WIDE
    exePacket[3]      = fab_chip.fabScalar.exePipe3.exePacket;
`endif
end
*/

/* Following maintains all the performance related counters. */
/*
always @(posedge clk)
begin: UPDATE_STATS
    int i;

    if (CYCLE_COUNT > 10)
    begin
        fetch1_stall      = fetch1_stall   + fab_chip.fabScalar.fs1.stall_i;
        ctiq_stall        = ctiq_stall     + fab_chip.fabScalar.fs2.ctiQueueFull;
        instBuf_stall     = instBuf_stall  + fab_chip.fabScalar.instBuf.instBufferFull;
        freelist_stall    = freelist_stall + fab_chip.fabScalar.rename.freeListEmpty;
        backend_stall     = backend_stall  + fab_chip.fabScalar.dispatch.stall;
        ldq_stall         = ldq_stall      + fab_chip.fabScalar.dispatch.loadStall;
        stq_stall         = stq_stall      + fab_chip.fabScalar.dispatch.storeStall;
        iq_stall          = iq_stall       + fab_chip.fabScalar.dispatch.iqStall;
        rob_stall         = rob_stall      + fab_chip.fabScalar.dispatch.alStall;

        btb_miss          = btb_miss       + (~fab_chip.fabScalar.fs1.stall_i & fab_chip.fabScalar.fs1.fs2RecoverFlag_i);
        btb_miss_rtn      = btb_miss_rtn   + (~fab_chip.fabScalar.fs1.stall_i &
                                               fab_chip.fabScalar.fs1.fs2MissedReturn_i &
                                               fab_chip.fabScalar.fs1.fs2RecoverFlag_i);
        for (i = 0; i < `COMMIT_WIDTH; i++)
        begin
            br_count        = br_count       + ((fab_chip.fabScalar.activeList.totalCommit >= (i+1)) & fab_chip.fabScalar.activeList.ctrlAl[i][5]);
            ld_count        = ld_count       + fab_chip.fabScalar.activeList.commitLoad_o[i];
        end

        br_mispredict_count =  br_mispredict_count + fab_chip.fabScalar.activeList.mispredFlag_reg;

        load_violation_count = load_violation_count + fab_chip.fabScalar.activeList.violateFlag_reg;

        ib_count  = ib_count  + fab_chip.fabScalar.instBuf.instCount;
        fl_count  = fl_count  + fab_chip.fabScalar.rename.specfreelist.freeListCnt;
        iq_count  = iq_count  + fab_chip.fabScalar.cntInstIssueQ;
        ldq_count = ldq_count + fab_chip.fabScalar.ldqCount;
        stq_count = stq_count + fab_chip.fabScalar.stqCount;
        al_count  = al_count  + fab_chip.fabScalar.activeListCnt;
        
        commit_1  = commit_1  + ((fab_chip.fabScalar.activeList.totalCommit == 1) ? 1'h1: 1'h0);
        commit_2  = commit_2  + ((fab_chip.fabScalar.activeList.totalCommit == 2) ? 1'h1: 1'h0);
        commit_3  = commit_3  + ((fab_chip.fabScalar.activeList.totalCommit == 3) ? 1'h1: 1'h0);
        commit_4  = commit_4  + ((fab_chip.fabScalar.activeList.totalCommit == 4) ? 1'h1: 1'h0);

    end
end
*/
always @(posedge clk)
begin: END_SIMULATION

    if (COMMIT_COUNT >= SIM_STOP_COUNT)
    begin

        ipc = $itor(COMMIT_COUNT)/$itor(CYCLE_COUNT);

/*
        // Before the simulator is terminated, print all the stats:
        $display(" Fetch1-Stall:%d \n Ctiq-Stall:%d \n InstBuff-Stall:%d \n FreeList-Stall:%d \n SMT-Stall:%d \n Backend-Stall:%d \n LDQ-Stall:%d \n STQ-Stall:%d \n IQ-Stall:%d \n ROB-Stall:%d\n",
        fetch1_stall,
        ctiq_stall,
        instBuf_stall,
        freelist_stall,
        smt_stall,
        backend_stall,
        ldq_stall,
        stq_stall,
        iq_stall,
        rob_stall);

        $display("stat_num_corr        %d", `stat_num_corr);
        $display("stat_num_pred        %d", `stat_num_pred);
        $display("stat_num_cond_corr   %d", `stat_num_cond_corr);
        $display("stat_num_cond_pred   %d", `stat_num_cond_pred);
        $display("stat_num_return_corr %d", `stat_num_return_corr);
        $display("stat_num_return_pred %d", `stat_num_return_pred);
        $display("");

        ib_avg    = ib_count/(CYCLE_COUNT-10.0);
        fl_avg    = fl_count/(CYCLE_COUNT-10.0);
        iq_avg    = iq_count/(CYCLE_COUNT-10.0);
        ldq_avg   = ldq_count/(CYCLE_COUNT-10.0);
        stq_avg   = stq_count/(CYCLE_COUNT-10.0);
        al_avg    = al_count/(CYCLE_COUNT-10.0);

        $write(" IB-avg: %2.1f\n", ib_avg); 
        $write(" FL-avg: %2.1f\n", fl_avg); 
        $write(" IQ-avg: %2.1f\n", iq_avg); 
        $write(" LDQ-avg: %2.1f\n", ldq_avg); 
        $write(" STQ-avg: %2.1f\n", stq_avg); 
        $write(" AL-avg: %2.1f\n", al_avg); 
      */
        $display("Cycle Count:%d Commit Count:%d    IPC:%2.2f     BTB-Miss:%d BTB-Miss-Rtn:%d  Br-Count:%d Br-Mispredict:%d Ld Count:%d Ld Violation:%d",
        CYCLE_COUNT,
        COMMIT_COUNT,
        ipc,
        btb_miss,
        btb_miss_rtn,
        br_count,
        br_mispredict_count,
        ld_count,
        load_violation_count);
      /*
        `ifdef DUMP_STATS
        ib_avg    = ib_count/(CYCLE_COUNT-10.0);
        fl_avg    = fl_count/(CYCLE_COUNT-10.0);
        iq_avg    = iq_count/(CYCLE_COUNT-10.0);
        ldq_avg   = ldq_count/(CYCLE_COUNT-10.0);
        stq_avg   = stq_count/(CYCLE_COUNT-10.0);
        al_avg    = al_count/(CYCLE_COUNT-10.0);

        $fwrite(fd16, "%d, ", CYCLE_COUNT); 
        $fwrite(fd16, "%d, ", COMMIT_COUNT); 

        $fwrite(fd16, "%2.3f, ", ib_avg); 
        $fwrite(fd16, "%2.3f, ", fl_avg); 
        $fwrite(fd16, "%2.3f, ", iq_avg); 
        $fwrite(fd16, "%2.4f, ", ldq_avg); 
        $fwrite(fd16, "%2.4f, ", stq_avg); 
        $fwrite(fd16, "%2.3f, ", al_avg); 

        $fwrite(fd16, "%d, ", fetch1_stall); 
        $fwrite(fd16, "%d, ", ctiq_stall); 
        $fwrite(fd16, "%d, ", instBuf_stall); 
        $fwrite(fd16, "%d, ", freelist_stall); 
        $fwrite(fd16, "%d, ", backend_stall); 
        $fwrite(fd16, "%d, ", ldq_stall); 
        $fwrite(fd16, "%d, ", stq_stall); 
        $fwrite(fd16, "%d, ", iq_stall); 
        $fwrite(fd16, "%d, ", rob_stall); 

        $fwrite(fd16, "%d, ", btb_miss); 
        $fwrite(fd16, "%d, ", btb_miss_rtn); 
        $fwrite(fd16, "%d, ", br_count); 
        $fwrite(fd16, "%d, ", br_mispredict_count); 
        $fwrite(fd16, "%d, ", load_violation_count); 

        $fwrite(fd16, "%d, ", `stat_num_corr);
        $fwrite(fd16, "%d, ", `stat_num_pred);
        $fwrite(fd16, "%d, ", `stat_num_cond_corr);
        $fwrite(fd16, "%d, ", `stat_num_cond_pred);
        $fwrite(fd16, "%d, ", `stat_num_return_corr);
        $fwrite(fd16, "%d, ", `stat_num_return_pred);

        $fwrite(fd16, "%d, ", commit_1); 
        $fwrite(fd16, "%d, ", commit_2); 
        $fwrite(fd16, "%d, ", commit_3); 
        $fwrite(fd16, "%d\n", commit_4); 
        `endif

        $fclose(fd0);
        $fclose(fd1);
        $fclose(fd2);
        $fclose(fd3);
        $fclose(fd4);
        $fclose(fd5);
        $fclose(fd6);
        $fclose(fd7);
        $fclose(fd8);
        $fclose(fd9);
        $fclose(fd10);
        $fclose(fd11);
        $fclose(fd12);
        $fclose(fd13);
        $fclose(fd14);
        $fclose(fd16);
        $fclose(fd17);
        $fclose(fd18);
        $fclose(fd19);
        $fclose(fd20);
        $fclose(fd21);
        $fclose(fd22);
        $fclose(fd23);

        //`endif
*/      
        $finish;
        read_AMT();
      `ifdef PERF_MON
        read_perf_mon();
      `endif  
    end
end

`ifdef PRINT_EN

/*  Prints top level related latches in a file every cycle. */
always @(posedge clk)
begin : FABSCALAR
    int i;

  if (PRINT)
  begin
        $fwrite(fd9, "------------------------------------------------------\n");
        $fwrite(fd9, "Cycle: %0d  Commit: %0d\n\n",CYCLE_COUNT, COMMIT_COUNT);

`ifdef DYNAMIC_CONFIG
        $fwrite(fd9, "stallFetch: %b\n\n", fab_chip.fabScalar.stallFetch);
`endif        

  end
end
`endif



`ifdef PRINT_EN
btbDataPkt                           btbData       [0:`FETCH_WIDTH-1];

always_comb
begin
    int i;
    for (i = 0; i < `FETCH_WIDTH; i++)
    begin
        btbData[i]  = fab_chip.fabScalar.fs1.btb.btbData[i];
    end
end

/*  Prints fetch1 stage related latches in a file every cycle. */
always @(posedge clk)
begin : FETCH1
    int i;

  if (PRINT)
  begin
        $fwrite(fd9, "------------------------------------------------------\n");
        $fwrite(fd9, "Cycle: %0d  Commit: %0d\n\n",CYCLE_COUNT, COMMIT_COUNT);

        $fwrite(fd9, "stall_i: %b\n\n", fab_chip.fabScalar.fs1.stall_i);

        $fwrite(fd9, "               -- Next PC --\n\n");
        
        $fwrite(fd9, "PC:             %08x\n",
                fab_chip.fabScalar.fs1.PC);

        $fwrite(fd9, "recoverPC_i:    %08x recoverFlag_i: %b mispredFlag_reg: %b violateFlag_reg: %b\n",
                fab_chip.fabScalar.fs1.recoverPC_i,
                fab_chip.fabScalar.fs1.recoverFlag_i,
                fab_chip.fabScalar.activeList.mispredFlag_reg,
                fab_chip.fabScalar.activeList.violateFlag_reg);

        $fwrite(fd9, "exceptionPC_i:  %08x exceptionFlag_i: %b\n",
                fab_chip.fabScalar.fs1.exceptionPC_i,
                fab_chip.fabScalar.fs1.exceptionFlag_i);

        $fwrite(fd9, "fs2RecoverPC_i: %08x fs2RecoverFlag_i: %b\n",
                fab_chip.fabScalar.fs1.fs2RecoverPC_i,
                fab_chip.fabScalar.fs1.fs2RecoverFlag_i);

        $fwrite(fd9, "nextPC:         %08x\n\n",
                fab_chip.fabScalar.fs1.nextPC);

        $fwrite(fd9, "takenVect:  %04b\n",
                fab_chip.fabScalar.fs1.takenVect);

        $fwrite(fd9, "addrRAS:    %08x\n\n",
                fab_chip.fabScalar.fs1.addrRAS);

        $fwrite(fd9, "               -- BTB --\n\n");
        
        $fwrite(fd9, "\nbtbData       ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd9, "     [%1d] ", i);

        $fwrite(fd9, "\ntag           ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd9, "%08x ", btbData[i].tag);

        $fwrite(fd9, "\ntakenPC       ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd9, "%08x ", btbData[i].takenPC);

        $fwrite(fd9, "\nctrlType      ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd9, "%08x ", btbData[i].ctrlType);

        $fwrite(fd9, "\nvalid         ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd9, "%08x ", btbData[i].valid);

        $fwrite(fd9, "\n\nupdatePC_i:     %08x\n",
                fab_chip.fabScalar.fs1.updatePC_i);

        $fwrite(fd9, "updateNPC_i:    %08x\n",
                fab_chip.fabScalar.fs1.updateNPC_i);

        $fwrite(fd9, "updateBrType_i: %x\n",
                fab_chip.fabScalar.fs1.updateBrType_i);

        $fwrite(fd9, "updateDir_i:    %b\n",
                fab_chip.fabScalar.fs1.updateDir_i);

        $fwrite(fd9, "updateEn_i:     %b\n\n",
                fab_chip.fabScalar.fs1.updateEn_i);


        $fwrite(fd9, "               -- BP --\n\n");
        
        $fwrite(fd9, "predDir:    %04b\n",
                fab_chip.fabScalar.fs1.predDir);

        $fwrite(fd9, "instOffset[0]:    %x\n",
                fab_chip.fabScalar.fs1.bp.instOffset[0]);

        $fwrite(fd9, "rdAddr         ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd9, "%x ", fab_chip.fabScalar.fs1.bp.rdAddr[i]);

        $fwrite(fd9, "\nrdData         ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd9, "%x ", fab_chip.fabScalar.fs1.bp.rdData[i]);

        $fwrite(fd9, "\npredCounter    ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd9, "%x ", fab_chip.fabScalar.fs1.bp.predCounter[i]);

        $fwrite(fd9, "\n\nwrAddr:        %x\n",
                fab_chip.fabScalar.fs1.bp.wrAddr);

        $fwrite(fd9, "\nwrData:        %x\n",
                fab_chip.fabScalar.fs1.bp.wrData);

        $fwrite(fd9, "\nwrEn         ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd9, "%x ", fab_chip.fabScalar.fs1.bp.wrEn[i]);


        $fwrite(fd9, "\n\n               -- RAS --\n\n");
        
        $fwrite(fd9, "pushAddr:   %08x\n",
                fab_chip.fabScalar.fs1.pushAddr);

        $fwrite(fd9, "pushRAS:   %b  popRAS: %b\n",
                fab_chip.fabScalar.fs1.pushRAS,
                fab_chip.fabScalar.fs1.popRAS);

        $fwrite(fd9, "\n\n");

        if (fab_chip.fabScalar.instBufferFull)
            $fwrite(fd9, "instBufferFull:%b\n",
                    fab_chip.fabScalar.instBufferFull);

    if (fab_chip.fabScalar.ctiQueueFull)
      $fwrite(fd9, "ctiQueueFull:%b\n",
              fab_chip.fabScalar.ctiQueueFull);

    if (fab_chip.fabScalar.fs1.recoverFlag_i)

    if(fab_chip.fabScalar.fs1.ras.pop_i)
      $fwrite(fd9, "BTB hit for Rtr instr, spec_tos:%d, Pop Addr: %x",
              fab_chip.fabScalar.fs1.ras.spec_tos,
              fab_chip.fabScalar.fs1.ras.addrRAS_o);

    if (fab_chip.fabScalar.fs1.ras.push_i)
      $fwrite(fd9, "BTB hit for CALL instr, Push Addr: %x",
              fab_chip.fabScalar.fs1.ras.pushAddr_i);

    $fwrite(fd9, "RAS POP Addr:%x\n",
            fab_chip.fabScalar.fs1.ras.addrRAS_o);

    if (fab_chip.fabScalar.fs1.fs2RecoverFlag_i)
      $fwrite(fd9, "Fetch-2 fix BTB miss (target addr): %h\n",
              fab_chip.fabScalar.fs1.fs2RecoverPC_i);

        $fwrite(fd9, "\n\n\n");
  end
end
`endif


`ifdef PRINT_EN
/* Prints fetch2/Ctrl Queue related latches in a file every cycle. */
always_ff @(posedge clk) 
begin : FETCH2
    int i;

  if (PRINT)
  begin
        $fwrite(fd14, "------------------------------------------------------\n");
        $fwrite(fd14, "Cycle: %0d  Commit: %0d\n\n\n",CYCLE_COUNT, COMMIT_COUNT);

    if (fab_chip.fabScalar.fs2.ctiQueue.stall_i)
    begin
      $fwrite(fd14, "Fetch2 is stalled ....\n");
    end

    if (fab_chip.fabScalar.fs2.ctiQueueFull_o)
    begin
      $fwrite(fd14, "CTI Queue is full ....\n");
    end

    $fwrite(fd14, "\n");

    $fwrite(fd14, "Control vector:%b fs1Ready:%b\n",
            fab_chip.fabScalar.fs2.ctiQueue.ctrlVect_i,
            fab_chip.fabScalar.fs2.ctiQueue.fs1Ready_i);


    $fwrite(fd14, "\n");

    $fwrite(fd14, "ctiq Tag0:%d ",
            fab_chip.fabScalar.fs2.ctiQueue.ctiID_o[0]);

`ifdef FETCH_TWO_WIDE
    $fwrite(fd14, "ctiq Tag1:%d ",
            fab_chip.fabScalar.fs2.ctiQueue.ctiID_o[1]);
`endif

`ifdef FETCH_THREE_WIDE
    $fwrite(fd14, "ctiq Tag2:%d ",
            fab_chip.fabScalar.fs2.ctiQueue.ctiID_o[2]);
`endif

`ifdef FETCH_FOUR_WIDE
    $fwrite(fd14, "ctiq Tag3:%d ",
            fab_chip.fabScalar.fs2.ctiQueue.ctiID_o[3]);
`endif

`ifdef FETCH_FIVE_WIDE
    $fwrite(fd14, "ctiq Tag4:%d ",
            fab_chip.fabScalar.fs2.ctiQueue.ctiID_o[4]);
`endif

`ifdef FETCH_SIX_WIDE
    $fwrite(fd14, "ctiq Tag5:%d ",
            fab_chip.fabScalar.fs2.ctiQueue.ctiID_o[5]);
`endif

`ifdef FETCH_SEVEN_WIDE
    $fwrite(fd14, "ctiq Tag6:%d ",
            fab_chip.fabScalar.fs2.ctiQueue.ctiID_o[6]);
`endif

`ifdef FETCH_EIGHT_WIDE
    $fwrite(fd14, "ctiq Tag7:%d ",
            fab_chip.fabScalar.fs2.ctiQueue.ctiID_o[7]);
`endif

        $fwrite(fd14, "\nupdateCounter_i:   %x\n",
                fab_chip.fabScalar.fs1.bp.updateCounter_i);

        $fwrite(fd14, "\ncti.headPtr:       %x\n",
                fab_chip.fabScalar.fs2.ctiQueue.headPtr);

        $fwrite(fd14, "\nctiq.ctiID            ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd14, "%x ", fab_chip.fabScalar.fs2.ctiQueue.ctiID[i]);

        $fwrite(fd14, "\nctiq.predCounter_i    ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd14, "%x ", fab_chip.fabScalar.fs2.ctiQueue.predCounter_i[i]);

        $fwrite(fd14, "\nctiq.ctrlVect_i       ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd14, "%x ", fab_chip.fabScalar.fs2.ctiQueue.ctrlVect_i[i]);

    $fwrite(fd14, "\n\n");

    if (fab_chip.fabScalar.fs2.ctiQueue.exeCtrlValid_i) begin
      $fwrite(fd14, "\nwriting back a control instruction.....\n");

      $fwrite(fd14,"ctiq index:%d target addr:%h br outcome:%b\n\n",
              fab_chip.fabScalar.fs2.ctiQueue.exeCtiID_i,
              fab_chip.fabScalar.fs2.ctiQueue.exeCtrlNPC_i,
              fab_chip.fabScalar.fs2.ctiQueue.exeCtrlDir_i);
    end

    if (fab_chip.fabScalar.fs2.ctiQueue.recoverFlag_i)
    begin
      $fwrite(fd14, "Recovery Flag is High....\n\n");
    end

    if (fab_chip.fabScalar.fs2.ctiQueue.updateEn_o)
    begin
      $fwrite(fd14, "\nupdating the BTB and BPB.....\n");

      $fwrite(fd14, "updatePC:%h updateNPC: %h updateCtrlType:%b updateDir:%b\n\n",
              fab_chip.fabScalar.fs2.ctiQueue.updatePC_o,
              fab_chip.fabScalar.fs2.ctiQueue.updateNPC_o,
              fab_chip.fabScalar.fs2.ctiQueue.updateCtrlType_o,
              fab_chip.fabScalar.fs2.updateDir_o);
    end

    $fwrite(fd14, "ctiq=> headptr:%d tailptr:%d commitPtr:%d instcount:%d commitCnt:%d\n",
            fab_chip.fabScalar.fs2.ctiQueue.headPtr,
            fab_chip.fabScalar.fs2.ctiQueue.tailPtr,
            fab_chip.fabScalar.fs2.ctiQueue.commitPtr,
            fab_chip.fabScalar.fs2.ctiQueue.ctrlCount,
            fab_chip.fabScalar.fs2.ctiQueue.commitCnt);

    $fwrite(fd14, "\n");
  end
end



/*  Prints decode stage related latches in a file every cycle. */
decPkt                     decPacket [0:`FETCH_WIDTH-1];
renPkt                     ibPacket [0:2*`FETCH_WIDTH-1];

always_comb
begin
    int i;
    for (i = 0; i < `FETCH_WIDTH; i++)
    begin
        decPacket[i]    = fab_chip.fabScalar.decPacket_l1[i];
        ibPacket[2*i]   = fab_chip.fabScalar.ibPacket[2*i];
        ibPacket[2*i+1] = fab_chip.fabScalar.ibPacket[2*i+1];
    end
end

always_ff @(posedge clk)
begin : DECODE
    int i;

    if (PRINT)
    begin
        $fwrite(fd2, "------------------------------------------------------\n");
        $fwrite(fd2, "Cycle: %0d  Commit: %0d\n\n\n",CYCLE_COUNT, COMMIT_COUNT);

        $fwrite(fd2, "fs2Ready_i: %b\n", fab_chip.fabScalar.decode.fs2Ready_i);

        $fwrite(fd2, "\n               -- decPackets --\n");
        
        $fwrite(fd2, "\ndecPacket_i   ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd2, "     [%1d] ", i);

        $fwrite(fd2, "\npc:           ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd2, "%08x ", decPacket[i].pc);

        $fwrite(fd2, "\nctrlType:     ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd2, "      %2x ", decPacket[i].ctrlType);

        $fwrite(fd2, "\nctiID:        ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd2, "      %2x ", decPacket[i].ctiID);

        $fwrite(fd2, "\npredNPC:      ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd2, "%08x ", decPacket[i].predNPC);

        $fwrite(fd2, "\npredDir:      ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd2, "       %1x ", decPacket[i].predDir);

        $fwrite(fd2, "\nvalid:        ");
        for (i = 0; i < `FETCH_WIDTH; i++)
            $fwrite(fd2, "       %1x ", decPacket[i].valid);


        $fwrite(fd2, "\n\n               -- ibPackets --\n");
        
        $fwrite(fd2, "\nibPacket_o    ");
        for (i = 0; i < 2*`FETCH_WIDTH; i++)
            $fwrite(fd2, "     [%1d] ", i);

        $fwrite(fd2, "\npc:           ");
        for (i = 0; i < 2*`FETCH_WIDTH; i++)
            $fwrite(fd2, "%08x ", ibPacket[i].pc);

        $fwrite(fd2, "\nopcode:       ");
        for (i = 0; i < 2*`FETCH_WIDTH; i++)
            $fwrite(fd2, "      %2x ",  ibPacket[i].opcode);

        $fwrite(fd2, "\nlogDest (V):  ");
        for (i = 0; i < 2*`FETCH_WIDTH; i++)
            $fwrite(fd2, "  %2x (%d) ", ibPacket[i].logDest, ibPacket[i].logDestValid);

        $fwrite(fd2, "\nlogSrc1 (V):  ");
        for (i = 0; i < 2*`FETCH_WIDTH; i++)
            $fwrite(fd2, "  %2x (%d) ", ibPacket[i].logSrc1, ibPacket[i].logSrc1Valid);

        $fwrite(fd2, "\nlogSrc2 (V):  ");
        for (i = 0; i < 2*`FETCH_WIDTH; i++)
            $fwrite(fd2, "  %2x (%d) ", ibPacket[i].logSrc2, ibPacket[i].logSrc2Valid);

        $fwrite(fd2, "\nimmed (V):    ");
        for (i = 0; i < 2*`FETCH_WIDTH; i++)
            $fwrite(fd2, "%04x (%d) ", ibPacket[i].immed, ibPacket[i].immedValid);

        $fwrite(fd2, "\nisLoad:       ");
        for (i = 0; i < 2*`FETCH_WIDTH; i++)
            $fwrite(fd2, "       %1x ", ibPacket[i].isLoad);

        $fwrite(fd2, "\nisStore:      ");
        for (i = 0; i < 2*`FETCH_WIDTH; i++)
            $fwrite(fd2, "       %1x ", ibPacket[i].isStore);

        $fwrite(fd2, "\nldstSize:     ");
        for (i = 0; i < 2*`FETCH_WIDTH; i++)
            $fwrite(fd2, "       %1x ", ibPacket[i].ldstSize);

        $fwrite(fd2, "\nctrlType:     ");
        for (i = 0; i < 2*`FETCH_WIDTH; i++)
            $fwrite(fd2, "      %2x ", ibPacket[i].ctrlType);

        $fwrite(fd2, "\nctiID:        ");
        for (i = 0; i < 2*`FETCH_WIDTH; i++)
            $fwrite(fd2, "      %2x ", ibPacket[i].ctiID);

        $fwrite(fd2, "\npredNPC:      ");
        for (i = 0; i < 2*`FETCH_WIDTH; i++)
            $fwrite(fd2, "%08x ", ibPacket[i].predNPC);

        $fwrite(fd2, "\npredDir:      ");
        for (i = 0; i < 2*`FETCH_WIDTH; i++)
            $fwrite(fd2, "       %1x ", ibPacket[i].predDir);

        $fwrite(fd2, "\nvalid:        ");
        for (i = 0; i < 2*`FETCH_WIDTH; i++)
            $fwrite(fd2, "       %1x ", ibPacket[i].valid);

        $fwrite(fd2, "\n\n\n");

    end
end


/*  Prints Instruction Buffer stage related latches in a file every cycle. */
always @(posedge clk)
begin:INSTBUF

  if (PRINT)
  begin
        $fwrite(fd1, "------------------------------------------------------\n");
        $fwrite(fd1, "Cycle: %0d  Commit: %0d\n\n\n",CYCLE_COUNT, COMMIT_COUNT);

    $fwrite(fd1, "Inst Buffer Full:%b freelistEmpty:%b stallFrontEnd:%b\n",
            fab_chip.fabScalar.instBuf.stallFetch_i,
            fab_chip.fabScalar.freeListEmpty,
            fab_chip.fabScalar.stallfrontEnd);

    $fwrite(fd1, "\n");

    $fwrite(fd1, "Decode Ready=%b\n",
            fab_chip.fabScalar.instBuf.decodeReady_i);

    $fwrite(fd1, "instbuffer head=%d instbuffer tail=%d inst count=%d\n",
            fab_chip.fabScalar.instBuf.headPtr,
            fab_chip.fabScalar.instBuf.tailPtr,
            fab_chip.fabScalar.instBuf.instCount);

    $fwrite(fd1, "instBufferReady_o:%b\n",
            fab_chip.fabScalar.instBuf.instBufferReady_o);

    if (fab_chip.fabScalar.recoverFlag)
      $fwrite(fd1, "recoverFlag_i is High\n");

    if (fab_chip.fabScalar.instBuf.flush_i)
      $fwrite(fd1, "flush_i is High\n");

    if (fab_chip.fabScalar.instBuf.instCount > `INST_QUEUE)
    begin
      $fwrite(fd1, "Instruction Buffer overflow\n");
      $display("\n** Cycle: %d Instruction Buffer Overflow **\n",CYCLE_COUNT);
    end

    $fwrite(fd1,"\n");
  end
end


/*  Prints rename stage related latches in a file every cycle. */
disPkt                     disPacket [0:`DISPATCH_WIDTH-1];
phys_reg                   freedPhyReg [0:`COMMIT_WIDTH-1];

always_comb
begin
    int i;
    for (i = 0; i < `DISPATCH_WIDTH; i++)
    begin
        disPacket[i]    = fab_chip.fabScalar.disPacket[i];
        freedPhyReg[i]  = fab_chip.fabScalar.rename.specfreelist.freedPhyReg_i[i];
    end
end

always @(posedge clk)
begin:RENAME
    int i;

  if (PRINT)
  begin
        $fwrite(fd0, "------------------------------------------------------\n");
        $fwrite(fd0, "Cycle: %0d  Commit: %0d\n\n\n",CYCLE_COUNT, COMMIT_COUNT);

        $fwrite(fd0, "Decode Ready: %b\n",
                fab_chip.fabScalar.rename.decodeReady_i);
                /* fab_chip.fabScalar.rename.branchCount_i); */

    $fwrite(fd0, "freeListEmpty: %b\n",
            fab_chip.fabScalar.rename.freeListEmpty);

        /* disPacket_o */
        $fwrite(fd0, "disPacket_o   ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd0, "     [%1d] ", i);

        $fwrite(fd0, "\npc:           ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd0, "%08x ", disPacket[i].pc);

        $fwrite(fd0, "\nopcode:       ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd0, "      %2x ",  disPacket[i].opcode);

        $fwrite(fd0, "\nfu:           ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd0, "       %1x ", disPacket[i].fu);

        $fwrite(fd0, "\nlogDest:      ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd0, "      %2x ", disPacket[i].logDest);

        $fwrite(fd0, "\nphyDest (V):  ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd0, "  %2x (%d) ", disPacket[i].phyDest, disPacket[i].phyDestValid);

        $fwrite(fd0, "\nphySrc1 (V):  ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd0, "  %2x (%d) ", disPacket[i].phySrc1, disPacket[i].phySrc1Valid);

        $fwrite(fd0, "\nphySrc2 (V):  ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd0, "  %2x (%d) ", disPacket[i].phySrc2, disPacket[i].phySrc2Valid);

        $fwrite(fd0, "\nimmed (V):    ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd0, "%04x (%d) ", disPacket[i].immed, disPacket[i].immedValid);

        $fwrite(fd0, "\nisLoad:       ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd0, "       %1x ", disPacket[i].isLoad);

        $fwrite(fd0, "\nisStore:      ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd0, "       %1x ", disPacket[i].isStore);

        $fwrite(fd0, "\nldstSize:     ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd0, "       %1x ", disPacket[i].ldstSize);

        $fwrite(fd0, "\nctiID:        ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd0, "      %2x ", disPacket[i].ctiID);

        $fwrite(fd0, "\npredNPC:      ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd0, "%08x ", disPacket[i].predNPC);

        $fwrite(fd0, "\npredDir:      ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd0, "       %1x ", disPacket[i].predDir);

        $fwrite(fd0, "\n\nrename ready:%b\n\n", fab_chip.fabScalar.rename.renameReady_o);

        $fwrite(fd0, "               -- Free List (Popped) --\n\n");

        $fwrite(fd0, "freeListHead: %x\n", fab_chip.fabScalar.rename.specfreelist.freeListHead);
        $fwrite(fd0, "freeListTail: %x\n", fab_chip.fabScalar.rename.specfreelist.freeListTail);
        $fwrite(fd0, "freeListCnt: d%d\n", fab_chip.fabScalar.rename.specfreelist.freeListCnt);
        $fwrite(fd0, "pushNumber: d%d\n", fab_chip.fabScalar.rename.specfreelist.pushNumber);
        
        $fwrite(fd0, "\nrdAddr:       ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd0, "      %2x ", fab_chip.fabScalar.rename.specfreelist.readAddr[i]);

        $fwrite(fd0, "\nfreePhyReg:   ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd0, "      %2x ", fab_chip.fabScalar.rename.specfreelist.freePhyReg[i]);

        $fwrite(fd0, "\n\n\n               -- Free List (Pushed) --\n\n");

        $fwrite(fd0, "\nfreedPhyReg (V): ");
        for (i = 0; i < `COMMIT_WIDTH; i++)
            $fwrite(fd0, "      %2x ", freedPhyReg[i].reg_id, freedPhyReg[i].valid);

    $fwrite(fd0,"\n\n\n");
  end
end
`endif


`ifdef PRINT_EN
/* Prints dispatch related signals and latch value. */
disPkt                           disPacket_l1 [0:`DISPATCH_WIDTH-1];
iqPkt                            iqPacket  [0:`DISPATCH_WIDTH-1];
alPkt                            alPacket  [0:`DISPATCH_WIDTH-1];
lsqPkt                           lsqPacket [0:`DISPATCH_WIDTH-1];

always_comb
begin
    int i;
    for (i = 0; i < `DISPATCH_WIDTH; i++)
    begin
        disPacket_l1[i]               = fab_chip.fabScalar.disPacket_l1[i];
        iqPacket[i]                = fab_chip.fabScalar.iqPacket[i];
        alPacket[i]                = fab_chip.fabScalar.alPacket[i];
        lsqPacket[i]               = fab_chip.fabScalar.lsqPacket[i];
    end
end

always_ff @(posedge clk)
begin:DISPATCH
    int i;

    if (PRINT)
    begin
        $fwrite(fd3, "----------------------------------------------------------------------\n");
        $fwrite(fd3, "Cycle: %d Commit Count: %d\n\n", CYCLE_COUNT, COMMIT_COUNT);

        /* disPacket_i */
        $fwrite(fd3, "disPacket_i   ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "     [%1d] ", i);

        $fwrite(fd3, "\npc:           ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "%08x ", disPacket_l1[i].pc);

        $fwrite(fd3, "\nopcode:       ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "      %2x ",  disPacket_l1[i].opcode);

        $fwrite(fd3, "\nfu:           ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "       %1x ", disPacket_l1[i].fu);

        $fwrite(fd3, "\nlogDest:      ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "      %2x ", disPacket_l1[i].logDest);

        $fwrite(fd3, "\nphyDest (V):  ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "  %2x (%d) ", disPacket_l1[i].phyDest, disPacket_l1[i].phyDestValid);

        $fwrite(fd3, "\nphySrc1 (V):  ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "  %2x (%d) ", disPacket_l1[i].phySrc1, disPacket_l1[i].phySrc1Valid);

        $fwrite(fd3, "\nphySrc2 (V):  ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "  %2x (%d) ", disPacket_l1[i].phySrc2, disPacket_l1[i].phySrc2Valid);

        $fwrite(fd3, "\nimmed (V):    ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "%04x (%d) ", disPacket_l1[i].immed, disPacket_l1[i].immedValid);

        $fwrite(fd3, "\nisLoad:       ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "       %1x ", disPacket_l1[i].isLoad);

        $fwrite(fd3, "\nisStore:      ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "       %1x ", disPacket_l1[i].isStore);

        $fwrite(fd3, "\nldstSize:     ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "       %1x ", disPacket_l1[i].ldstSize);

        $fwrite(fd3, "\nctiID:        ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "      %2x ", disPacket_l1[i].ctiID);

        $fwrite(fd3, "\npredNPC:      ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "%08x ", disPacket_l1[i].predNPC);

        $fwrite(fd3, "\npredDir:      ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "       %1x ", disPacket_l1[i].predDir);

        /* iqPacket_o */
        $fwrite(fd3, "\n\niqPacket_o    ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "     [%1d] ", i);

        $fwrite(fd3, "\npc:           ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "%08x ", iqPacket[i].pc);

        $fwrite(fd3, "\nopcode:       ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "      %2x ",  iqPacket[i].opcode);

        $fwrite(fd3, "\nfu:           ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "       %1x ", iqPacket[i].fu);

        $fwrite(fd3, "\nphyDest (V):  ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "  %2x (%d) ", iqPacket[i].phyDest, iqPacket[i].phyDestValid);

        $fwrite(fd3, "\nphySrc1 (V):  ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "  %2x (%d) ", iqPacket[i].phySrc1, iqPacket[i].phySrc1Valid);

        $fwrite(fd3, "\nphySrc2 (V):  ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "  %2x (%d) ", iqPacket[i].phySrc2, iqPacket[i].phySrc2Valid);

        $fwrite(fd3, "\nimmed (V):    ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "%04x (%d) ", iqPacket[i].immed, iqPacket[i].immedValid);

        $fwrite(fd3, "\nisLoad:       ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "       %1x ", iqPacket[i].isLoad);

        $fwrite(fd3, "\nisStore:      ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "       %1x ", iqPacket[i].isStore);

        $fwrite(fd3, "\nldstSize:     ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "       %1x ", iqPacket[i].ldstSize);

        $fwrite(fd3, "\nctiID:        ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "      %2x ", iqPacket[i].ctiID);

        $fwrite(fd3, "\npredNPC:      ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "%08x ", iqPacket[i].predNPC);

        $fwrite(fd3, "\npredDir:      ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd3, "       %1x ", iqPacket[i].predDir);


    $fwrite(fd3, "\n\nloadCnt: d%d storeCnt: d%d\n",
            fab_chip.fabScalar.dispatch.loadCnt,
            fab_chip.fabScalar.dispatch.storeCnt);

    $fwrite(fd3, "backendReady_o: %b\n",
            fab_chip.fabScalar.dispatch.backEndReady_o);

    if (fab_chip.fabScalar.dispatch.loadStall)       $fwrite(fd3,"LDQ Stall\n");
    if (fab_chip.fabScalar.dispatch.storeStall)      $fwrite(fd3,"STQ Stall\n");
    if (fab_chip.fabScalar.dispatch.iqStall)         $fwrite(fd3,"IQ Stall: IQ Cnt:%d\n",
                                                    fab_chip.fabScalar.dispatch.issueQueueCnt_i);
    if (fab_chip.fabScalar.dispatch.alStall)         $fwrite(fd3,"Active List Stall\n");
    if (~fab_chip.fabScalar.dispatch.renameReady_i)  $fwrite(fd3,"renameReady_i Stall\n");


`ifdef ENABLE_LD_VIOLATION_PRED
    $fwrite(fd3, "predictLdViolation: %b\n",
            fab_chip.fabScalar.dispatch.predLoadVio);

    if (fab_chip.fabScalar.dispatch.ldVioPred.loadViolation_i && fab_chip.fabScalar.dispatch.ldVioPred.recoverFlag_i)
    begin
      $fwrite(fd3, "Update Load Violation Predictor\n");

      $fwrite(fd3, "PC:0x%x Addr:0x%x Tag:0x%x\n",
              fab_chip.fabScalar.dispatch.ldVioPred.recoverPC_i,
              fab_chip.fabScalar.dispatch.ldVioPred.predAddr0wr,
              fab_chip.fabScalar.dispatch.ldVioPred.predTag0wr);
    end
`endif
    $fwrite(fd3,"\n",);
  end
end
`endif


`ifdef PRINT_EN
phys_reg                        phyDest  [0:`DISPATCH_WIDTH-1];
iqEntryPkt                      iqFreeEntry [0:`DISPATCH_WIDTH-1];

iqEntryPkt                      iqFreedEntry   [0:`ISSUE_WIDTH-1];
iqEntryPkt                      iqGrantedEntry [0:`ISSUE_WIDTH-1];
payloadPkt                      rrPacket       [0:`ISSUE_WIDTH-1];

always_comb
begin
    int i;
    for (i = 0; i < `DISPATCH_WIDTH; i++)
    begin
        phyDest[i]     = fab_chip.fabScalar.phyDest[i];
        iqFreeEntry[i] = fab_chip.fabScalar.issueq.freeEntry[i];
    end

    for (i = 0; i < `ISSUE_WIDTH; i++)
    begin
        iqFreedEntry[i] = fab_chip.fabScalar.issueq.freedEntry[i];
        iqGrantedEntry[i] = fab_chip.fabScalar.issueq.grantedEntry[i];
        rrPacket[i]     = fab_chip.fabScalar.rrPacket[i];
    end
end

/* Prints issue queue related signals and latch values. */
always_ff @(posedge clk)
begin: ISSUEQ
  int i;

    if (PRINT)
    begin
        $fwrite(fd5, "------------------------------------------------------\n");
        $fwrite(fd5, "Cycle: %0d  Commit: %0d\n\n\n",CYCLE_COUNT, COMMIT_COUNT);

`ifdef DYNAMIC_CONFIG
        $fwrite(fd7, "dispatchLaneActive_i: %x\n",
        fab_chip.fabScalar.issueq.dispatchLaneActive_i);

        $fwrite(fd7, "issueLaneActive_i: %x\n",
        fab_chip.fabScalar.issueq.issueLaneActive_i);
`endif        

        $fwrite(fd5, "               -- Dispatched Instructions --\n\n");
        
        $fwrite(fd5, "backEndReady_i:          %b\n", fab_chip.fabScalar.issueq.backEndReady_i);

        /* iqPacket_i */
        $fwrite(fd5, "iqPacket_i        ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "     [%1d] ", i);

        $fwrite(fd5, "\npc:               ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "%08x ", iqPacket[i].pc);

        $fwrite(fd5, "\nopcode:           ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "      %2x ",  iqPacket[i].opcode);

        $fwrite(fd5, "\nfu:               ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "       %1x ", iqPacket[i].fu);

        $fwrite(fd5, "\nphyDest (V):      ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "  %2x (%d) ", iqPacket[i].phyDest, iqPacket[i].phyDestValid);

        $fwrite(fd5, "\nphySrc1 (V):      ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "  %2x (%d) ", iqPacket[i].phySrc1, iqPacket[i].phySrc1Valid);

        $fwrite(fd5, "\nphySrc2 (V):      ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "  %2x (%d) ", iqPacket[i].phySrc2, iqPacket[i].phySrc2Valid);

        $fwrite(fd5, "\nimmed (V):        ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "%04x (%d) ", iqPacket[i].immed, iqPacket[i].immedValid);

        $fwrite(fd5, "\nisLoad:           ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "       %1x ", iqPacket[i].isLoad);

        $fwrite(fd5, "\nisStore:          ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "       %1x ", iqPacket[i].isStore);

        $fwrite(fd5, "\nldstSize:         ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "       %1x ", iqPacket[i].ldstSize);

        $fwrite(fd5, "\nctiID:            ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "      %2x ", iqPacket[i].ctiID);

        $fwrite(fd5, "\npredNPC:          ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "%08x ", iqPacket[i].predNPC);

        $fwrite(fd5, "\npredDir:          ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "       %1x ", iqPacket[i].predDir);

        $fwrite(fd5, "\nfreeEntry:        ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "     d%2d ", iqFreeEntry[i].id);

        $fwrite(fd5, "\nlsqID:            ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "      %2x ", fab_chip.fabScalar.lsqID[i]);

        $fwrite(fd5, "\nalID:             ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "      %2x ", fab_chip.fabScalar.alID[i]);

        /* phyDest_i */
        $fwrite(fd5, "\n\nphyDest_i         ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "     [%1d] ", i);

        $fwrite(fd5, "\nreg_id (V):       ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "  %2x (%1x) ", phyDest[i].reg_id, phyDest[i].valid);

        $fwrite(fd5, "\nnewSrc1Ready:     ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "       %b ", fab_chip.fabScalar.issueq.newSrc1Ready[i]);
 
        $fwrite(fd5, "\nnewSrc2Ready:     ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd5, "       %b ", fab_chip.fabScalar.issueq.newSrc2Ready[i]);

        $fwrite(fd5, "\nrsrTag:        ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
        begin
            $fwrite(fd5, "       %b ",fab_chip.fabScalar.issueq.rsrTag[i]);
        end 

        $fwrite(fd5, "\nrsrTag_t:    ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
        begin
            `ifndef DYNAMIC_CONFIG
              $fwrite(fd5, "       %b ",fab_chip.fabScalar.issueq.rsr.rsrTag_o[i]);
            `else
            `endif
        end
 
        $fwrite(fd5, "\nISsimple_t:    ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
        begin
            $fwrite(fd5, "       %b ",fab_chip.fabScalar.issueq.ISsimple_t[i]);
        end


        /* IQ Freelist */

        $fwrite(fd5, "\n\n               -- IQ Freelist --\n\n");

        $fwrite(fd5, "issueQCount: d%d headPtr: d%d tailPtr: d%d\n",
                fab_chip.fabScalar.issueq.issueQfreelist.issueQCount,
                fab_chip.fabScalar.issueq.issueQfreelist.headPtr,
                fab_chip.fabScalar.issueq.issueQfreelist.tailPtr);


        /* Wakeup */

        $fwrite(fd5, "\n\n               -- Wakeup --\n\n");

        $fwrite(fd5, "phyRegValidVect: %b\n\n", fab_chip.fabScalar.issueq.phyRegValidVect);
        
        $fwrite(fd5, "rsrTag (V):      ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
        begin
            $fwrite(fd5, "%2x (%b) ",
                    fab_chip.fabScalar.issueq.rsrTag[i][`SIZE_PHYSICAL_LOG:1],
                    fab_chip.fabScalar.issueq.rsrTag[i][0]);
        end

        //$fwrite(fd5, "\n\niqValidVect:     %b\n", fab_chip.fabScalar.issueq.iqValidVect);
        $fwrite(fd5, "src1MatchVect:   %b\n",     fab_chip.fabScalar.issueq.src1MatchVect);
        //$fwrite(fd5, "src1Valid_t1:    %b\n",     fab_chip.fabScalar.issueq.src1Valid_t1);
        //$fwrite(fd5, "src1ValidVect:   %b\n",     fab_chip.fabScalar.issueq.src1ValidVect);

        //$fwrite(fd5, "\n\niqValidVect:     %b\n", fab_chip.fabScalar.issueq.iqValidVect);
        $fwrite(fd5, "src2MatchVect:   %b\n",     fab_chip.fabScalar.issueq.src2MatchVect);
        //$fwrite(fd5, "src2Valid_t1:    %b\n",     fab_chip.fabScalar.issueq.src2Valid_t1);
        //$fwrite(fd5, "src2ValidVect:   %b\n",     fab_chip.fabScalar.issueq.src2ValidVect);


        /* Select */

        $fwrite(fd5, "\n\n               -- Select --\n\n");

        //$fwrite(fd5, "iqValidVect:     %b\n", fab_chip.fabScalar.issueq.iqValidVect);
        //$fwrite(fd5, "src1ValidVect:   %b\n", fab_chip.fabScalar.issueq.src1ValidVect);
        //$fwrite(fd5, "src2ValidVect:   %b\n", fab_chip.fabScalar.issueq.src2ValidVect);
        $fwrite(fd5, "reqVect:         %b\n", fab_chip.fabScalar.issueq.reqVect);
        `ifndef DYNAMIC_CONFIG
          $fwrite(fd5, "reqVectFU0:      %b\n", fab_chip.fabScalar.issueq.reqVectFU0);
          $fwrite(fd5, "reqVectFU1:      %b\n", fab_chip.fabScalar.issueq.reqVectFU1);
          $fwrite(fd5, "reqVectFU2:      %b\n", fab_chip.fabScalar.issueq.reqVectFU2);
          `ifdef ISSUE_FOUR_WIDE
            $fwrite(fd5, "reqVectFU3:      %b\n", fab_chip.fabScalar.issueq.reqVectFU3);
          `endif
          `ifdef ISSUE_FIVE_WIDE
            $fwrite(fd5, "reqVectFU4:      %b\n", fab_chip.fabScalar.issueq.reqVectFU4);
          `endif
        `else
        `endif

        //$fwrite(fd5, "grantedVect:     %b\n", fab_chip.fabScalar.issueq.grantedVect);

        /* rrPacket_o */
        $fwrite(fd5, "\nrrPacket_o        ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd5, "     [%1d] ", i);

        $fwrite(fd5, "\npc:               ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd5, "%08x ", rrPacket[i].pc);

        $fwrite(fd5, "\nopcode:           ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd5, "      %2x ",  rrPacket[i].opcode);

        $fwrite(fd5, "\nphyDest:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd5, "      %2x ", rrPacket[i].phyDest);

        $fwrite(fd5, "\nphySrc1:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd5, "      %2x ", rrPacket[i].phySrc1);

        $fwrite(fd5, "\nphySrc2:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd5, "      %2x ", rrPacket[i].phySrc2);

        $fwrite(fd5, "\nimmed:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd5, "    %04x ", rrPacket[i].immed);

        $fwrite(fd5, "\nlsqID:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd5, "      %2x ", rrPacket[i].lsqID);

        $fwrite(fd5, "\nalID:             ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd5, "      %2x ", rrPacket[i].alID);

        $fwrite(fd5, "\nldstSize:         ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd5, "       %1x ", rrPacket[i].ldstSize);

        $fwrite(fd5, "\nctiID:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd5, "      %2x ", rrPacket[i].ctiID);

        $fwrite(fd5, "\npredNPC:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd5, "%08x ", rrPacket[i].predNPC);

        $fwrite(fd5, "\npredDir:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd5, "       %1x ", rrPacket[i].predDir);

        $fwrite(fd5, "\ngrantedEntry (V): ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd5, "  %2x (%1d) ", iqGrantedEntry[i].id, iqGrantedEntry[i].valid);

        $fwrite(fd5,"\n\n");

        //$fwrite(fd5, "freedVect:       %b\n", fab_chip.fabScalar.issueq.freedVect);
        $fwrite(fd5, "freedEntry (V): ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd5, "  %2x (%1d) ", iqFreedEntry[i].id, iqFreedEntry[i].valid);
        
        $fwrite(fd5,"\n");
        /* for (i = 0;i< `NO_OF_COMPLEX; i++) */
        /* $fwrite(fd5,"issue_simple[%x] : %b    ",i,fab_chip.fabScalar.issueq.issue_simple[i]); */    
/*
        $fwrite(fd5,"\n\n");
        $fwrite(fd5,"RSR1 (V) :");
        for (i = 0;i < `FU1_LATENCY;i++)
            $fwrite(fd5,"   %2x (%1d) ",fab_chip.fabScalar.issueq.rsr.RSR_CALU1[i],fab_chip.fabScalar.issueq.rsr.RSR_CALU_VALID1[i]);
        $fwrite(fd5,"\n\n");
        
        $fwrite(fd5,"RSR2 (V) :");
        for (i = 0;i < `FU1_LATENCY;i++)
            $fwrite(fd5,"   %2x (%1d) ",fab_chip.fabScalar.issueq.rsr.RSR_CALU2[i],fab_chip.fabScalar.issueq.rsr.RSR_CALU_VALID2[i]);
*/
        $fwrite(fd5,"\n\n\n");
    end
end
`endif /* PRINT_EN */


`ifdef PRINT_EN
payloadPkt                      rrPacket_l1    [0:`ISSUE_WIDTH-1];
bypassPkt                       bypassPacket   [0:`ISSUE_WIDTH-1];
/* fuPkt                           exePacket      [0:`ISSUE_WIDTH-1]; */

always_comb
begin
    int i;
    for (i = 0; i < `ISSUE_WIDTH; i++)
    begin
        rrPacket_l1[i]  = fab_chip.fabScalar.rrPacket_l1[i];
        bypassPacket[i] = fab_chip.fabScalar.bypassPacket[i];
    end
end

/* Prints register read related signals and latch value. */
always_ff @(posedge clk)
begin : REG_READ
    int i;

    if (PRINT)
    begin

        $fwrite(fd6, "------------------------------------------------------\n");
        $fwrite(fd6, "Cycle: %0d  Commit: %0d\n\n",CYCLE_COUNT, COMMIT_COUNT);

        $fwrite(fd6, "               -- rrPacket_i --\n");

        /* rrPacket_i */
        $fwrite(fd6, "\nrrPacket_i        ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "     [%1d] ", i);

        $fwrite(fd6, "\npc:               ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "%08x ", rrPacket_l1[i].pc);

        $fwrite(fd6, "\nopcode:           ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "      %2x ",  rrPacket_l1[i].opcode);

        $fwrite(fd6, "\nphyDest:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "      %2x ", rrPacket_l1[i].phyDest);

        $fwrite(fd6, "\nphySrc1:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "      %2x ", rrPacket_l1[i].phySrc1);

        $fwrite(fd6, "\nphySrc2:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "      %2x ", rrPacket_l1[i].phySrc2);

        $fwrite(fd6, "\nimmed:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "    %04x ", rrPacket_l1[i].immed);

        $fwrite(fd6, "\nlsqID:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "      %2x ", rrPacket_l1[i].lsqID);

        $fwrite(fd6, "\nalID:             ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "      %2x ", rrPacket_l1[i].alID);

        /* $fwrite(fd6, "\nldstSize:         "); */
        /* for (i = 0; i < `ISSUE_WIDTH; i++) */
        /*     $fwrite(fd6, "       %1x ", rrPacket_l1[i].ldstSize); */

        $fwrite(fd6, "\nctiID:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "      %2x ", rrPacket_l1[i].ctiID);

        $fwrite(fd6, "\npredNPC:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "%08x ", rrPacket_l1[i].predNPC);

        $fwrite(fd6, "\npredDir:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "       %1x ", rrPacket_l1[i].predDir);

        $fwrite(fd6, "\nvalid:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "       %1x ", rrPacket_l1[i].valid);


        $fwrite(fd6, "\n\n               -- bypassPacket_i --\n");

        /* rrPacket_i */
        $fwrite(fd6, "\nbypassPacket_i    ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "     [%1d] ", i);

        $fwrite(fd6, "\ntag:              ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "      %2x ", bypassPacket[i].tag);

        $fwrite(fd6, "\ndata:             ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "%08x ",  bypassPacket[i].data);

        $fwrite(fd6, "\nvalid:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "       %1x ", bypassPacket[i].valid);


        $fwrite(fd6, "\n\n               -- exePacket_o --\n");

        /* rrPacket_i */
        $fwrite(fd6, "\nexePacket_o       ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "     [%1d] ", i);

        $fwrite(fd6, "\npc:               ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "%08x ", exePacket[i].pc);

        $fwrite(fd6, "\nopcode:           ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "      %2x ",  exePacket[i].opcode);

        $fwrite(fd6, "\nphyDest:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "      %2x ", exePacket[i].phyDest);

        $fwrite(fd6, "\nphySrc1:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "      %2x ", exePacket[i].phySrc1);

        $fwrite(fd6, "\nsrc1Data:         ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "%08x ", exePacket[i].src1Data);

        $fwrite(fd6, "\nphySrc2:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "      %2x ", exePacket[i].phySrc2);

        $fwrite(fd6, "\nsrc2Data:         ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "%08x ", exePacket[i].src2Data);

        $fwrite(fd6, "\nimmed:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "    %04x ", exePacket[i].immed);

        $fwrite(fd6, "\nlsqID:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "      %2x ", exePacket[i].lsqID);

        $fwrite(fd6, "\nalID:             ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "      %2x ", exePacket[i].alID);

        /* $fwrite(fd6, "\nldstSize:         "); */
        /* for (i = 0; i < `ISSUE_WIDTH; i++) */
        /*     $fwrite(fd6, "       %1x ", exePacket[i].ldstSize); */

        $fwrite(fd6, "\nctiID:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "      %2x ", exePacket[i].ctiID);

        $fwrite(fd6, "\npredNPC:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "%08x ", exePacket[i].predNPC);

        $fwrite(fd6, "\npredDir:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "       %1x ", exePacket[i].predDir);

        $fwrite(fd6, "\nvalid:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd6, "       %1x ", exePacket[i].valid);

        $fwrite(fd6, "\n\n\n");

    end
end
`endif // PRINT_EN


`ifdef PRINT_EN
reg  [`SIZE_PHYSICAL_LOG-1:0]               src1Addr_byte0 [0:`ISSUE_WIDTH-1];
reg  [`SIZE_PHYSICAL_LOG-1:0]               src1Addr_byte1 [0:`ISSUE_WIDTH-1];
reg  [`SIZE_PHYSICAL_LOG-1:0]               src1Addr_byte2 [0:`ISSUE_WIDTH-1];
reg  [`SIZE_PHYSICAL_LOG-1:0]               src1Addr_byte3 [0:`ISSUE_WIDTH-1];
reg  [`SIZE_PHYSICAL_LOG-1:0]               src2Addr_byte0 [0:`ISSUE_WIDTH-1];
reg  [`SIZE_PHYSICAL_LOG-1:0]               src2Addr_byte1 [0:`ISSUE_WIDTH-1];
reg  [`SIZE_PHYSICAL_LOG-1:0]               src2Addr_byte2 [0:`ISSUE_WIDTH-1];
reg  [`SIZE_PHYSICAL_LOG-1:0]               src2Addr_byte3 [0:`ISSUE_WIDTH-1];
reg  [`SIZE_PHYSICAL_LOG-1:0]               destAddr_byte0 [0:`ISSUE_WIDTH-1];
reg  [`SIZE_PHYSICAL_LOG-1:0]               destAddr_byte1 [0:`ISSUE_WIDTH-1];
reg  [`SIZE_PHYSICAL_LOG-1:0]               destAddr_byte2 [0:`ISSUE_WIDTH-1];
reg  [`SIZE_PHYSICAL_LOG-1:0]               destAddr_byte3 [0:`ISSUE_WIDTH-1];

always_comb
begin
    int i, j;
    for (i = 0; i < `ISSUE_WIDTH; i++)
    begin
        for (j = 0; j < `SIZE_PHYSICAL_TABLE; j++)
        begin
            if (fab_chip.fabScalar.registerfile.src1Addr_byte0[i][j])
            begin
                src1Addr_byte0[i]              = j;
            end

            if (fab_chip.fabScalar.registerfile.src1Addr_byte1[i][j])
            begin
                src1Addr_byte1[i]              = j;
            end

            if (fab_chip.fabScalar.registerfile.src1Addr_byte2[i][j])
            begin
                src1Addr_byte2[i]              = j;
            end

            if (fab_chip.fabScalar.registerfile.src1Addr_byte3[i][j])
            begin
                src1Addr_byte3[i]              = j;
            end


            if (fab_chip.fabScalar.registerfile.src2Addr_byte0[i][j])
            begin
                src2Addr_byte0[i]              = j;
            end

            if (fab_chip.fabScalar.registerfile.src2Addr_byte1[i][j])
            begin
                src2Addr_byte1[i]              = j;
            end

            if (fab_chip.fabScalar.registerfile.src2Addr_byte2[i][j])
            begin
                src2Addr_byte2[i]              = j;
            end

            if (fab_chip.fabScalar.registerfile.src2Addr_byte3[i][j])
            begin
                src2Addr_byte3[i]              = j;
            end


            if (fab_chip.fabScalar.registerfile.destAddr_byte0[i][j])
            begin
                destAddr_byte0[i]              = j;
            end

            if (fab_chip.fabScalar.registerfile.destAddr_byte1[i][j])
            begin
                destAddr_byte1[i]              = j;
            end

            if (fab_chip.fabScalar.registerfile.destAddr_byte2[i][j])
            begin
                destAddr_byte2[i]              = j;
            end

            if (fab_chip.fabScalar.registerfile.destAddr_byte3[i][j])
            begin
                destAddr_byte3[i]              = j;
            end
        end
    end
end


/* Prints register read related signals and latch value. */
always_ff @(posedge clk)
begin : PHY_REG_FILE
    int i;

    if (PRINT)
    begin

        $fwrite(fd23, "------------------------------------------------------\n");
        $fwrite(fd23, "Cycle: %0d  Commit: %0d\n\n",CYCLE_COUNT, COMMIT_COUNT);

        $fwrite(fd23, "               -- Read --\n");

        /* Read */
        $fwrite(fd23, "\n                  ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "     [%1d] ", i);

        $fwrite(fd23, "\nsrc1Addr_byte0:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", src1Addr_byte0[i]);

        $fwrite(fd23, "\nsrc1Data_byte0:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", fab_chip.fabScalar.registerfile.src1Data_byte0_o[i]);

        $fwrite(fd23, "\n\nsrc1Addr_byte1:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", src1Addr_byte1[i]);

        $fwrite(fd23, "\nsrc1Data_byte1:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", fab_chip.fabScalar.registerfile.src1Data_byte1_o[i]);

        $fwrite(fd23, "\n\nsrc1Addr_byte2:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", src1Addr_byte2[i]);

        $fwrite(fd23, "\nsrc1Data_byte2:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", fab_chip.fabScalar.registerfile.src1Data_byte2_o[i]);

        $fwrite(fd23, "\n\nsrc1Addr_byte3:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", src1Addr_byte3[i]);

        $fwrite(fd23, "\nsrc1Data_byte3:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", fab_chip.fabScalar.registerfile.src1Data_byte3_o[i]);


        $fwrite(fd23, "\n\nsrc2Addr_byte0:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", src2Addr_byte0[i]);

        $fwrite(fd23, "\nsrc2Data_byte0:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", fab_chip.fabScalar.registerfile.src2Data_byte0_o[i]);

        $fwrite(fd23, "\n\nsrc2Addr_byte1:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", src2Addr_byte1[i]);

        $fwrite(fd23, "\nsrc2Data_byte1:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", fab_chip.fabScalar.registerfile.src2Data_byte1_o[i]);

        $fwrite(fd23, "\n\nsrc2Addr_byte2:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", src2Addr_byte2[i]);

        $fwrite(fd23, "\nsrc2Data_byte2:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", fab_chip.fabScalar.registerfile.src2Data_byte2_o[i]);

        $fwrite(fd23, "\n\nsrc2Addr_byte3:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", src2Addr_byte3[i]);

        $fwrite(fd23, "\nsrc2Data_byte3:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", fab_chip.fabScalar.registerfile.src2Data_byte3_o[i]);

        $fwrite(fd23, "\n\n\n               -- Write --\n");

        /* Write */
        $fwrite(fd23, "\n                  ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "     [%1d] ", i);

        $fwrite(fd23, "\ndestAddr_byte0:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", destAddr_byte0[i]);

        $fwrite(fd23, "\ndestData_byte0:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", fab_chip.fabScalar.registerfile.destData_byte0[i]);

        $fwrite(fd23, "\ndestWe_byte0:     ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "       %1x ", fab_chip.fabScalar.registerfile.destWe_byte0[i]);

        $fwrite(fd23, "\n\ndestAddr_byte1:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", destAddr_byte1[i]);

        $fwrite(fd23, "\ndestData_byte1:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", fab_chip.fabScalar.registerfile.destData_byte1[i]);

        $fwrite(fd23, "\ndestWe_byte1:     ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "       %1x ", fab_chip.fabScalar.registerfile.destWe_byte1[i]);

        $fwrite(fd23, "\n\ndestAddr_byte2:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", destAddr_byte2[i]);

        $fwrite(fd23, "\ndestData_byte2:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", fab_chip.fabScalar.registerfile.destData_byte2[i]);

        $fwrite(fd23, "\ndestWe_byte2:     ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "       %1x ", fab_chip.fabScalar.registerfile.destWe_byte2[i]);

        $fwrite(fd23, "\n\ndestAddr_byte3:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", destAddr_byte3[i]);

        $fwrite(fd23, "\ndestData_byte3:   ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "      %02x ", fab_chip.fabScalar.registerfile.destData_byte3[i]);

        $fwrite(fd23, "\ndestWe_byte3:     ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd23, "       %1x ", fab_chip.fabScalar.registerfile.destWe_byte3[i]);

        $fwrite(fd23, "\n\n\n");

    end
end
`endif // PRINT_EN


`ifdef PRINT_EN
/* Prints functional units */
fuPkt                           exePacket_l1   [0:`ISSUE_WIDTH-1];
wbPkt                           wbPacket       [0:`ISSUE_WIDTH-1];
reg  [31:0]                     src1Data       [0:`ISSUE_WIDTH-1];
reg  [31:0]                     src2Data       [0:`ISSUE_WIDTH-1];

always_comb
begin
    int i;

    exePacket_l1[0]   = fab_chip.fabScalar.exePipe0.exePacket_l1;
    wbPacket[0]       = fab_chip.fabScalar.wbPacket;
    src1Data[0]       = fab_chip.fabScalar.exePipe0.execute.src1Data;
    src2Data[0]       = fab_chip.fabScalar.exePipe0.execute.src2Data;

    exePacket_l1[1]   = fab_chip.fabScalar.exePipe1.exePacket_l1;
    wbPacket[1]       = fab_chip.fabScalar.exePipe1.wbPacket;
    src1Data[1]       = fab_chip.fabScalar.exePipe1.execute.src1Data;
    src2Data[1]       = fab_chip.fabScalar.exePipe1.execute.src2Data;

    exePacket_l1[2]   = fab_chip.fabScalar.exePipe2.exePacket_l1;
    wbPacket[2]       = fab_chip.fabScalar.exePipe2.wbPacket;
    src1Data[2]       = fab_chip.fabScalar.exePipe2.execute.src1Data;
    src2Data[2]       = fab_chip.fabScalar.exePipe2.execute.src2Data;


`ifdef ISSUE_FOUR_WIDE
    exePacket_l1[3]   = fab_chip.fabScalar.exePipe3.exePacket_l1;
    wbPacket[3]       = fab_chip.fabScalar.exePipe3.wbPacket;
    src1Data[3]       = fab_chip.fabScalar.exePipe3.execute.src1Data;
    src2Data[3]       = fab_chip.fabScalar.exePipe3.execute.src2Data;
`endif

`ifdef ISSUE_FIVE_WIDE
    exePacket_l1[4]   = fab_chip.fabScalar.exePipe4.exePacket_l1;
    wbPacket[4]       = fab_chip.fabScalar.exePipe4.wbPacket;
    src1Data[4]       = fab_chip.fabScalar.exePipe4.execute.src1Data;
    src2Data[4]       = fab_chip.fabScalar.exePipe4.execute.src2Data;
`endif

`ifdef ISSUE_SIX_WIDE
    exePacket_l1[5]   = fab_chip.fabScalar.exePipe5.exePacket_l1;
    wbPacket[5]       = fab_chip.fabScalar.exePipe5.wbPacket;
    src1Data[5]       = fab_chip.fabScalar.exePipe5.execute.src1Data;
    src2Data[5]       = fab_chip.fabScalar.exePipe5.execute.src2Data;
`endif

`ifdef ISSUE_SEVEN_WIDE
    exePacket_l1[6]   = fab_chip.fabScalar.exePipe6.exePacket_l1;
    wbPacket[6]       = fab_chip.fabScalar.exePipe6.wbPacket;
    src1Data[6]       = fab_chip.fabScalar.exePipe6.execute.src1Data;
    src2Data[6]       = fab_chip.fabScalar.exePipe6.execute.src2Data;
`endif

end


always_ff @(posedge clk)
begin : EXE
    int i;

    if (PRINT)
    begin

        $fwrite(fd13, "------------------------------------------------------\n");
        $fwrite(fd13, "Cycle: %0d  Commit: %0d\n\n", CYCLE_COUNT, COMMIT_COUNT);


        $fwrite(fd13, "               -- exePacket_i --\n");

        /* exePacket_l1_i */
        $fwrite(fd13, "\nexePacket_i       ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "     [%1d] ", i);

        $fwrite(fd13, "\npc:               ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "%08x ", exePacket_l1[i].pc);

        $fwrite(fd13, "\nopcode:           ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "      %2x ",  exePacket_l1[i].opcode);

        $fwrite(fd13, "\nphyDest:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "      %2x ", exePacket_l1[i].phyDest);

        $fwrite(fd13, "\nphySrc1:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "      %2x ", exePacket_l1[i].phySrc1);

        $fwrite(fd13, "\nsrc1Data:         ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "%08x ", exePacket_l1[i].src1Data);

        $fwrite(fd13, "\nphySrc2:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "      %2x ", exePacket_l1[i].phySrc2);

        $fwrite(fd13, "\nsrc2Data:         ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "%08x ", exePacket_l1[i].src2Data);

        $fwrite(fd13, "\nimmed:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "    %04x ", exePacket_l1[i].immed);

        $fwrite(fd13, "\nlsqID:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "      %2x ", exePacket_l1[i].lsqID);

        $fwrite(fd13, "\nalID:             ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "      %2x ", exePacket_l1[i].alID);

        $fwrite(fd13, "\nctiID:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "      %2x ", exePacket_l1[i].ctiID);

        $fwrite(fd13, "\npredNPC:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "%08x ", exePacket_l1[i].predNPC);

        $fwrite(fd13, "\npredDir:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "       %1x ", exePacket_l1[i].predDir);

        $fwrite(fd13, "\nvalid:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "       %1x ", exePacket_l1[i].valid);


        $fwrite(fd13, "\n\n               -- bypassPacket_i --\n");

        /* rrPacket_i */
        $fwrite(fd13, "\nbypassPacket_i    ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "     [%1d] ", i);

        $fwrite(fd13, "\ntag:              ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "      %2x ", bypassPacket[i].tag);

        $fwrite(fd13, "\ndata:             ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "%8x ",  bypassPacket[i].data);

        $fwrite(fd13, "\nvalid:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "       %1x ", bypassPacket[i].valid);


        $fwrite(fd13, "\n\nsrc1Data:         ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "%08x ", src1Data[i]);

        $fwrite(fd13, "\nsrc2Data:         ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "%08x ", src2Data[i]);


        $fwrite(fd13, "\n\n               -- wbPacket_o --\n");

        /* wbPacket_i */
        $fwrite(fd13, "\nwbPacket_i        ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "     [%1d] ", i);

        $fwrite(fd13, "\npc:               ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "%08x ", wbPacket[i].pc);

        $fwrite(fd13, "\nflags:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "      %2x ",  wbPacket[i].flags);

        $fwrite(fd13, "\nphyDest:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "      %2x ", wbPacket[i].phyDest);

        $fwrite(fd13, "\ndestData:         ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "%08x ", wbPacket[i].destData);

        $fwrite(fd13, "\nalID:             ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "      %2x ", wbPacket[i].alID);

        $fwrite(fd13, "\nnextPC:           ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "%08x ", wbPacket[i].nextPC);

        $fwrite(fd13, "\nctrlType:         ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "      %2x ", wbPacket[i].ctrlType);

        $fwrite(fd13, "\nctrlDir:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "       %x ", wbPacket[i].ctrlDir);

        $fwrite(fd13, "\nctiID:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "      %2x ", wbPacket[i].ctiID);

        $fwrite(fd13, "\npredDir:          ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "       %1x ", wbPacket[i].predDir);

        $fwrite(fd13, "\nvalid:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd13, "       %1x ", wbPacket[i].valid);

        $fwrite(fd13, "\n\n\n");

    end
end
`endif // PRINT_EN


`ifdef PRINT_EN
/* Prints load-store related signals and latch value. */

memPkt                         memPacket;
memPkt                         replayPacket;

wbPkt                          lsuWbPacket;
ldVioPkt                       ldVioPacket;

always_comb
begin
    memPacket      = fab_chip.fabScalar.memPacket;
    replayPacket   = fab_chip.fabScalar.lsu.datapath.replayPacket;
    lsuWbPacket    = fab_chip.fabScalar.wbPacket;
    ldVioPacket    = fab_chip.fabScalar.ldVioPacket;
end


always @(posedge clk)
begin:LSU
    reg [`SIZE_LSQ_LOG-1:0]               lastMatch;
  reg [2+`SIZE_PC+`SIZE_RMT_LOG+2*`SIZE_PHYSICAL_LOG:0] val;
  int i;

  if (PRINT)
  begin
        $fwrite(fd10, "------------------------------------------------------\n");
        $fwrite(fd10, "Cycle: %0d  Commit: %0d\n\n\n",CYCLE_COUNT, COMMIT_COUNT);

        $fwrite(fd10, "               -- Dispatched Instructions --\n\n");
        
        $fwrite(fd10, "ldqHead_i:      %x\n", fab_chip.fabScalar.lsu.datapath.stx_path.ldqHead_i);
        $fwrite(fd10, "ldqTail_i:      %x\n", fab_chip.fabScalar.lsu.datapath.stx_path.ldqTail_i);
        $fwrite(fd10, "stqHead_i:      %x\n", fab_chip.fabScalar.lsu.datapath.ldx_path.stqHead_i);
        $fwrite(fd10, "stqTail_i:      %x\n", fab_chip.fabScalar.lsu.datapath.ldx_path.stqTail_i);
        $fwrite(fd10, "backEndReady_i: %b\n", fab_chip.fabScalar.lsu.backEndReady_i);
        $fwrite(fd10, "recoverFlag_i : %b\n", fab_chip.fabScalar.lsu.recoverFlag_i);

        /* lsqPacket_i */
        $fwrite(fd10, "lsqPacket_i       ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd10, "     [%1d] ", i);

        $fwrite(fd10, "\npredLoadVio:      ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd10, "       %1x ", lsqPacket[i].predLoadVio);

        $fwrite(fd10, "\nisLoad:           ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd10, "       %1x ", lsqPacket[i].isLoad);

        $fwrite(fd10, "\nisStore:          ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd10, "       %1x ", lsqPacket[i].isStore);

        $fwrite(fd10, "\nlsqID:            ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd10, "      %2x ", fab_chip.fabScalar.lsqID[i]);

        $fwrite(fd10, "\nldqID:            ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd10, "      %2x ", fab_chip.fabScalar.lsu.ldqID[i]);

        $fwrite(fd10, "\nstqID:            ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd10, "      %2x ", fab_chip.fabScalar.lsu.stqID[i]);

        $fwrite(fd10, "\nnextLd:            ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd10, "      %x ", fab_chip.fabScalar.lsu.datapath.nextLdIndex_i[i]);

        $fwrite(fd10, "\nlastSt:            ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd10, "      %x ", fab_chip.fabScalar.lsu.datapath.lastStIndex_i[i]);

        $fwrite(fd10, "\n\n\n               -- Executed Instructions --\n\n");
        
        /* memPacket_i */
        $fwrite(fd10, "memPacket_i       ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "     [%1d] ", i);

        $fwrite(fd10, "\nPC:            ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "      %x  ", memPacket.pc);

        $fwrite(fd10, "\nflags:            ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "      %2x ", memPacket.flags);

        $fwrite(fd10, "\nldstSize:         ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "       %1x ", memPacket.ldstSize);

        $fwrite(fd10, "\nphyDest:          ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "      %2x ", memPacket.phyDest);

        $fwrite(fd10, "\naddress:          ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "%08x ",     memPacket.address);

        $fwrite(fd10, "\nsrc2Data:         ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "%08x ",     memPacket.src2Data);

        $fwrite(fd10, "\nlsqID:            ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "      %2x ", memPacket.lsqID);

        $fwrite(fd10, "\nalID:             ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "      %2x ", memPacket.alID);

        $fwrite(fd10, "\nvalid:            ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "       %1x ", memPacket.valid);

        /* replayPacket_i */
        $fwrite(fd10, "\n\nreplayPacket       ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "     [%1d] ", i);

        $fwrite(fd10, "\nPC:            ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "      %x  ", replayPacket.pc);

        $fwrite(fd10, "\nflags:            ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "      %2x ", replayPacket.flags);

        $fwrite(fd10, "\nldstSize:         ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "       %1x ", replayPacket.ldstSize);

        $fwrite(fd10, "\nphyDest:          ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "      %2x ", replayPacket.phyDest);

        $fwrite(fd10, "\naddress:          ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "%08x ",     replayPacket.address);

        $fwrite(fd10, "\nsrc2Data:         ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "%08x ",     replayPacket.src2Data);

        $fwrite(fd10, "\nlsqID:            ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "      %2x ", replayPacket.lsqID);

        $fwrite(fd10, "\nalID:             ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "      %2x ", replayPacket.alID);

        $fwrite(fd10, "\nvalid:            ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "       %1x ", replayPacket.valid);

        $fwrite(fd10, "\n\n\nlastSt:            ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "       %x ", fab_chip.fabScalar.lsu.datapath.ldx_path.LD_DISAMBIGUATION.lastSt);


        /* lsuWbPacket_o */
        $fwrite(fd10, "\n\nlsuWbPacket_o        ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "     [%1d] ", i);

        $fwrite(fd10, "\npc:               ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "%08x ", lsuWbPacket.pc);

        $fwrite(fd10, "\nflags:            ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "      %2x ", lsuWbPacket.flags);

        $fwrite(fd10, "\nphyDest:          ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "      %2x ", lsuWbPacket.phyDest);

        $fwrite(fd10, "\ndestData:         ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "%08x ",     lsuWbPacket.destData);

        $fwrite(fd10, "\nalID:             ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "      %2x ", lsuWbPacket.alID);

        $fwrite(fd10, "\nvalid:            ");
        for (i = 0; i < 1; i++)
            $fwrite(fd10, "       %1x ", lsuWbPacket.valid);


        $fwrite(fd10, "\n\n\n               -- LD Disambiguation (LDX) --\n\n");

        $fwrite(fd10, "stqCount_i:  %x\n",
                fab_chip.fabScalar.lsu.datapath.ldx_path.stqCount_i);

        $fwrite(fd10, "stqAddrValid:  %b\n",
                fab_chip.fabScalar.lsu.datapath.ldx_path.stqAddrValid);

        $fwrite(fd10, "stqValid:  %b\n",
                fab_chip.fabScalar.lsu.control.stqValid);

        $fwrite(fd10, "vulnerableStVector_t1:  %b\n",
                fab_chip.fabScalar.lsu.datapath.ldx_path.LD_DISAMBIGUATION.vulnerableStVector_t1);

        $fwrite(fd10, "vulnerableStVector_t2:  %b\n",
                fab_chip.fabScalar.lsu.datapath.ldx_path.LD_DISAMBIGUATION.vulnerableStVector_t2);

        $fwrite(fd10, "vulnerableStVector:     %b\n",
                fab_chip.fabScalar.lsu.datapath.ldx_path.LD_DISAMBIGUATION.vulnerableStVector);

`ifndef DYNAMIC_CONFIG                
        $fwrite(fd10, "addr1MatchVector:       %b\n",
                fab_chip.fabScalar.lsu.datapath.ldx_path.LD_DISAMBIGUATION.addr1MatchVector);

        $fwrite(fd10, "addr2MatchVector:       %b\n",
                fab_chip.fabScalar.lsu.datapath.ldx_path.LD_DISAMBIGUATION.addr2MatchVector);
`else                
        $fwrite(fd10, "addr1MatchVector:       %b\n",
                fab_chip.fabScalar.lsu.datapath.ldx_path.addr1MatchVector);

        $fwrite(fd10, "addr2MatchVector:       %b\n",
                fab_chip.fabScalar.lsu.datapath.ldx_path.addr2MatchVector);
`endif

        $fwrite(fd10, "sizeMismatchVector:     %b\n",
                fab_chip.fabScalar.lsu.datapath.ldx_path.LD_DISAMBIGUATION.sizeMismatchVector);

        $fwrite(fd10, "forwardVector1:         %b\n",
                fab_chip.fabScalar.lsu.datapath.ldx_path.LD_DISAMBIGUATION.forwardVector1);

        $fwrite(fd10, "forwardVector2:         %b\n\n",
                fab_chip.fabScalar.lsu.datapath.ldx_path.LD_DISAMBIGUATION.forwardVector2);


`ifndef DYNAMIC_CONFIG        
        lastMatch = fab_chip.fabScalar.lsu.datapath.ldx_path.LD_DISAMBIGUATION.lastMatch;
`else
        lastMatch = fab_chip.fabScalar.lsu.datapath.ldx_path.lastMatch;
`endif
        $fwrite(fd10, "stqHit:         %b\n", fab_chip.fabScalar.lsu.datapath.ldx_path.stqHit);
        $fwrite(fd10, "lastMatch:      %x\n", lastMatch);
        $fwrite(fd10, "partialStMatch: %b\n", fab_chip.fabScalar.lsu.datapath.ldx_path.partialStMatch);
        $fwrite(fd10, "disambigStall:  %b\n\n", fab_chip.fabScalar.lsu.datapath.ldx_path.LD_DISAMBIGUATION.disambigStall);

        $fwrite(fd10, "loadDataValid_o: %b\n", fab_chip.fabScalar.lsu.datapath.ldx_path.loadDataValid_o);
        $fwrite(fd10, "dcacheData:  %08x\n", fab_chip.fabScalar.lsu.datapath.ldx_path.dcacheData);
`ifndef DYNAMIC_CONFIG        
        $fwrite(fd10, "stqData[%d]: %08x\n", lastMatch, fab_chip.fabScalar.lsu.datapath.ldx_path.stqData[lastMatch]);
`else        
        $fwrite(fd10, "stqData[%d]: %08x\n", lastMatch, fab_chip.fabScalar.lsu.datapath.ldx_path.stqHitData);
`endif
        $fwrite(fd10, "loadData_t:  %08x\n", fab_chip.fabScalar.lsu.datapath.ldx_path.loadData_t);
        $fwrite(fd10, "loadData_o:  %08x\n", fab_chip.fabScalar.lsu.datapath.ldx_path.loadData_o);
        

        $fwrite(fd10, "\n\n\n               -- LD Violation (STX) --\n\n");

        $fwrite(fd10, "ldqAddrValid:           %b\n",
                fab_chip.fabScalar.lsu.datapath.stx_path.ldqAddrValid);

        $fwrite(fd10, "ldqWriteBack:           %b\n",
                fab_chip.fabScalar.lsu.datapath.stx_path.ldqWriteBack);

        $fwrite(fd10, "vulnerableLdVector_t1:  %b\n",
                fab_chip.fabScalar.lsu.datapath.stx_path.LD_VIOLATION.vulnerableLdVector_t1);

        $fwrite(fd10, "vulnerableLdVector_t2:  %b\n",
                fab_chip.fabScalar.lsu.datapath.stx_path.LD_VIOLATION.vulnerableLdVector_t2);

        $fwrite(fd10, "vulnerableLdVector_t3:  %b\n",
                fab_chip.fabScalar.lsu.datapath.stx_path.LD_VIOLATION.vulnerableLdVector_t3);

        $fwrite(fd10, "vulnerableLdVector_t4:  %b\n",
                fab_chip.fabScalar.lsu.datapath.stx_path.LD_VIOLATION.vulnerableLdVector_t4);

        $fwrite(fd10, "matchVector_st:         %b\n",
                fab_chip.fabScalar.lsu.datapath.stx_path.LD_VIOLATION.matchVector_st);

`ifndef DYNAMIC_CONFIG
        $fwrite(fd10, "matchVector_st1:        %b\n",
                fab_chip.fabScalar.lsu.datapath.stx_path.LD_VIOLATION.matchVector_st1);
`else                
        $fwrite(fd10, "matchVector_st1:        %b\n",
                fab_chip.fabScalar.lsu.datapath.stx_path.matchVector_st1);
`endif

        $fwrite(fd10, "matchVector_st2:        %b\n",
                fab_chip.fabScalar.lsu.datapath.stx_path.LD_VIOLATION.matchVector_st2);

        $fwrite(fd10, "matchVector_st3:        %b\n",
                fab_chip.fabScalar.lsu.datapath.stx_path.LD_VIOLATION.matchVector_st3);

        $fwrite(fd10, "violateVector:          %b\n",
                fab_chip.fabScalar.lsu.datapath.stx_path.LD_VIOLATION.violateVector);


        $fwrite(fd10, "nextLoad:       %x\n", fab_chip.fabScalar.lsu.datapath.stx_path.LD_VIOLATION.nextLoad);
`ifndef DYNAMIC_CONFIG
        $fwrite(fd10, "firstMatch:     %x\n", fab_chip.fabScalar.lsu.datapath.stx_path.LD_VIOLATION.firstMatch);
`else                
        $fwrite(fd10, "firstMatch:     %x\n", fab_chip.fabScalar.lsu.datapath.stx_path.firstMatch);
`endif
        $fwrite(fd10, "agenLdqMatch:   %b\n", fab_chip.fabScalar.lsu.datapath.stx_path.LD_VIOLATION.agenLdqMatch);
        $fwrite(fd10, "violateLdValid: %x\n", fab_chip.fabScalar.lsu.datapath.stx_path.violateLdValid);
        $fwrite(fd10, "violateLdALid:  %x\n", fab_chip.fabScalar.lsu.datapath.stx_path.violateLdALid);
        
        $fwrite(fd10, "\n\n\n               -- Committed Instructions --\n\n");
        
        $fwrite(fd10, "stqHead_i:   %d\n", fab_chip.fabScalar.lsu.datapath.ldx_path.stqHead_i);
        $fwrite(fd10, "commitSt_i:  %x\n", fab_chip.fabScalar.lsu.datapath.ldx_path.commitSt_i);
        $fwrite(fd10, "stCommitAddr:  %x\n", fab_chip.fabScalar.lsu.datapath.ldx_path.stCommitAddr);
        $fwrite(fd10, "stCommitData:  %x\n", fab_chip.fabScalar.lsu.datapath.ldx_path.stCommitData);
        $fwrite(fd10, "commitStCount:  %x", fab_chip.fabScalar.lsu.control.commitStCount);
        $fwrite(fd10, "commitStIndex: ");
        for (i = 0; i < 4; i++)
        begin
          $fwrite(fd10, "  %x", fab_chip.fabScalar.lsu.control.commitStIndex[i]);
        end

        for (i = 0; i < `SIZE_LSQ; i++)
        begin
`ifndef DYNAMIC_CONFIG          
            $fwrite(fd10, "stqAddr[%0d]: %08x\n", i, {fab_chip.fabScalar.lsu.datapath.ldx_path.stqAddr1[i],
                                                      fab_chip.fabScalar.lsu.datapath.ldx_path.stqAddr2[i]});
`endif                                                      
        end
        
        for (i = 0; i < `SIZE_LSQ; i++)
        begin
`ifndef DYNAMIC_CONFIG          
            $fwrite(fd10, "stqData[%0d]: %08x\n", i, fab_chip.fabScalar.lsu.datapath.ldx_path.stqData[i]);
`endif
        end

    $fwrite(fd10, "commitLoad_i:  %b\n",
              fab_chip.fabScalar.lsu.commitLoad_i);

    $fwrite(fd10, "commitStore_i: %b\n",
              fab_chip.fabScalar.lsu.commitStore_i);

    $fwrite(fd10,"\n\n");
  end
end
`endif // 0



`ifdef PRINT_EN
ctrlPkt                         ctrlPacket [0:`ISSUE_WIDTH-1];
commitPkt                       amtPacket [0:`COMMIT_WIDTH-1];

always_comb
begin
    int i;
    for (i = 0; i < `ISSUE_WIDTH; i++)
    begin
        ctrlPacket[i]   = fab_chip.fabScalar.ctrlPacket[i];
    end

    for (i = 0; i < `COMMIT_WIDTH; i++)
    begin
        amtPacket[i]   = fab_chip.fabScalar.amtPacket[i];
    end
end

always_ff @(posedge clk)
begin: ACTIVE_LIST
    int i;

    if (PRINT)
    begin
        $fwrite(fd7, "------------------------------------------------------\n");
        $fwrite(fd7, "Cycle: %0d  Commit: %0d\n\n\n",CYCLE_COUNT, COMMIT_COUNT);

`ifdef DYNAMIC_CONFIG
        $fwrite(fd7, "dispatchLaneActive_i: %x\n",
        fab_chip.fabScalar.activeList.dispatchLaneActive_i);

        $fwrite(fd7, "issueLaneActive_i: %x\n",
        fab_chip.fabScalar.activeList.issueLaneActive_i);
`endif        

        $fwrite(fd7, "totalCommit: d%d\n",
        fab_chip.fabScalar.activeList.totalCommit);

        $fwrite(fd7, "alCount: d%d\n",
        fab_chip.fabScalar.activeList.alCount);

        $fwrite(fd7, "headPtr: %x tailPtr: %x\n",
        fab_chip.fabScalar.activeList.headPtr,
        fab_chip.fabScalar.activeList.tailPtr);

        $fwrite(fd7, "backEndReady_i: %b\n\n",
        fab_chip.fabScalar.activeList.backEndReady_i);

        $fwrite(fd7, "               -- Dispatched Instructions --\n\n");
        
        /* alPacket_i */
        $fwrite(fd7, "\nalPacket_i    ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd7, "     [%1d] ", i);

        $fwrite(fd7, "\npc:           ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd7, "%08x ", alPacket[i].pc);

        $fwrite(fd7, "\nlogDest:      ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd7, "      %2x ", alPacket[i].logDest);

        $fwrite(fd7, "\nphyDest (V):  ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd7, "  %2x (%d) ", alPacket[i].phyDest, alPacket[i].phyDestValid);

        $fwrite(fd7, "\nisLoad:       ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd7, "       %1x ", alPacket[i].isLoad);

        $fwrite(fd7, "\nisStore:      ");
        for (i = 0; i < `DISPATCH_WIDTH; i++)
            $fwrite(fd7, "       %1x ", alPacket[i].isStore);

        $fwrite(fd7, "\n\n\n               -- Executed Instructions --\n");

        $fwrite(fd7, "\nctrlPacket_i      ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd7, "     [%1d] ", i);

        $fwrite(fd7, "\nnextPC:           ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd7, "%08x ", ctrlPacket[i].nextPC);

        $fwrite(fd7, "\nalID:             ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd7, "      %2x ", ctrlPacket[i].alID);

        $fwrite(fd7, "\nflags:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd7, "      %2x ", ctrlPacket[i].flags);

        $fwrite(fd7, "\nvalid:            ");
        for (i = 0; i < `ISSUE_WIDTH; i++)
            $fwrite(fd7, "       %1x ", ctrlPacket[i].valid);
        
        
        $fwrite(fd7, "\n\n\n               -- Committing Instructions --\n\n");
        
        $fwrite(fd7, "              ");
        for (i = 0; i < `COMMIT_WIDTH; i++)
            $fwrite(fd7, "     [%1d] ", i);

        $fwrite(fd7, "\nmispredFlag:  "); 
        for (i = 0; i < `COMMIT_WIDTH; i++)
            $fwrite(fd7, "       %b ", fab_chip.fabScalar.activeList.mispredFlag[i]);

        $fwrite(fd7, "\nviolateFlag:  ");
        for (i = 0; i < `COMMIT_WIDTH; i++)
            $fwrite(fd7, "       %b ", fab_chip.fabScalar.activeList.violateFlag[i]);
        
        $fwrite(fd7, "\nexceptionFlag:");
        for (i = 0; i < `COMMIT_WIDTH; i++)
            $fwrite(fd7, "       %b ", fab_chip.fabScalar.activeList.exceptionFlag[i]);

        $fwrite(fd7, "\n\ncommitReady:  ");
        for (i = 0; i < `COMMIT_WIDTH; i++)
            $fwrite(fd7, "       %b ", fab_chip.fabScalar.activeList.commitReady[i]);

        $fwrite(fd7, "\ncommitVector: ");
        for (i = 0; i < `COMMIT_WIDTH; i++)
            $fwrite(fd7, "       %b ", fab_chip.fabScalar.activeList.commitVector[i]);


        $fwrite(fd7, "\n\namtPacket_o   ");
        for (i = 0; i < `COMMIT_WIDTH; i++)
            $fwrite(fd7, "     [%1d] ", i);

        $fwrite(fd7, "\nlogDest:      ");
        for (i = 0; i < `COMMIT_WIDTH; i++)
            $fwrite(fd7, "      %2x ", amtPacket[i].logDest);

        $fwrite(fd7, "\nphyDest:      ");
        for (i = 0; i < `COMMIT_WIDTH; i++)
            $fwrite(fd7, "      %2x ", amtPacket[i].phyDest);

        $fwrite(fd7, "\nvalid:        ");
        for (i = 0; i < `COMMIT_WIDTH; i++)
            $fwrite(fd7, "       %1x ", amtPacket[i].valid);

        $fwrite(fd7, "\npc:           ");
        for (i = 0; i < `COMMIT_WIDTH; i++)
            $fwrite(fd7, "%08x ", fab_chip.fabScalar.activeList.commitPC[i]);

        $fwrite(fd7, "\n\ncommitStore:  ");
        for (i = 0; i < `COMMIT_WIDTH; i++)
            $fwrite(fd7, "       %1x ", fab_chip.fabScalar.activeList.commitStore_o[i]);

        $fwrite(fd7, "\ncommitLoad:   ");
        for (i = 0; i < `COMMIT_WIDTH; i++)
            $fwrite(fd7, "       %1x ", fab_chip.fabScalar.activeList.commitLoad_o[i]);

        $fwrite(fd7, "\ncommitCti:    ");
        for (i = 0; i < `COMMIT_WIDTH; i++)
            $fwrite(fd7, "       %1x ", fab_chip.fabScalar.activeList.commitCti_o[i]);

        $fwrite(fd7,"\n\n");

        
        if (fab_chip.fabScalar.activeList.violateFlag_reg)
        begin
            $fwrite(fd7, "violateFlag_reg: %d recoverPC_o: %h\n",
            fab_chip.fabScalar.activeList.violateFlag_reg,
            fab_chip.fabScalar.activeList.recoverPC_o);
        end

        if (fab_chip.fabScalar.activeList.mispredFlag_reg)
        begin
            $fwrite(fd7,"mispredFlag_reg: %d recoverPC_o: %h\n",
            fab_chip.fabScalar.activeList.mispredFlag_reg,
            fab_chip.fabScalar.activeList.recoverPC_o);
        end

        if (fab_chip.fabScalar.activeList.exceptionFlag_reg)
        begin
            $fwrite(fd7,"exceptionFlag_reg: %d exceptionPC_o: %h\n",
            fab_chip.fabScalar.activeList.exceptionFlag_reg,
            fab_chip.fabScalar.activeList.exceptionPC_o);
        end

        $fwrite(fd7,"\n");
    end
end

`endif


`ifdef PNR_SIM

      fs2Pkt  [0:`FETCH_WIDTH-1]                   fs2Packet;
      fs2Pkt  [0:`FETCH_WIDTH-1]                   fs2Packet_l1;
      
      assign        fs2Packet     = fab_chip.any.fabScalar.fs1fs2.fs2Packet_i;
      assign        fs2Packet_l1  = fab_chip.any.fabScalar.fs1fs2.fs2Packet_o;
      
      decPkt  [0:`FETCH_WIDTH-1]                   decPacket;
      decPkt  [0:`FETCH_WIDTH-1]                   decPacket_l1;
      renPkt  [0:2*`FETCH_WIDTH-1]                 ibPacket;
      
      assign        decPacket     = fab_chip.any.fabScalar.fs2dec.decPacket_i;
      assign        decPacket_l1  = fab_chip.any.fabScalar.fs2dec.decPacket_o;
      assign        ibPacket      = fab_chip.any.fabScalar.decode.ibPacket_o;
      
      renPkt  [0:`DISPATCH_WIDTH-1]                renPacket;
      renPkt  [0:`DISPATCH_WIDTH-1]                renPacket_l1;
      
      assign        renPacket     = fab_chip.any.fabScalar.instBufRen.renPacket_i;
      assign        renPacket_l1  = fab_chip.any.fabScalar.instBufRen.renPacket_o;
      
      
      disPkt  [0:`DISPATCH_WIDTH-1]                     disPacket_l1;
      iqPkt   [0:`DISPATCH_WIDTH-1]                     iqPacket;
      alPkt   [0:`DISPATCH_WIDTH-1]                     alPacket;
      lsqPkt  [0:`DISPATCH_WIDTH-1]                     lsqPacket;
      
      assign        disPacket_l1                = fab_chip.any.fabScalar.renDis.disPacket_o;
      assign        iqPacket                    = fab_chip.any.fabScalar.dispatch.iqPacket_o;
      assign        alPacket                    = fab_chip.any.fabScalar.dispatch.alPacket_o;
      assign        lsqPacket                   = fab_chip.any.fabScalar.lsu.lsqPacket_i;
      
      iqEntryPkt    [0:`ISSUE_WIDTH-1]              iqGrantedEntry;
      iqEntryPkt    [0:`ISSUE_WIDTH-1]              iqFreedEntry  ;
      iqEntryPkt    [0:`DISPATCH_WIDTH-1]           iqFreeEntry   ;
      
      assign        iqGrantedEntry                = fab_chip.any.fabScalar.issueq.issueQfreelist.grantedEntry_i;
      assign        iqFreedEntry                  = fab_chip.any.fabScalar.issueq.issueQfreelist.freedEntry_o;
      assign        iqFreeEntry                   = fab_chip.any.fabScalar.issueq.issueQfreelist.freeEntry_o;
      
      payloadPkt                                    iqPldWrPacket [0:`DISPATCH_WIDTH-1];
        assign        iqPldWrPacket[0] = fab_chip.any.fabScalar.issueq.payloadRAM.data0wr_i;
      `ifdef DISPATCH_TWO_WIDE
        assign        iqPldWrPacket[1] = fab_chip.any.fabScalar.issueq.payloadRAM.data1wr_i;
      `endif
      `ifdef DISPATCH_THREE_WIDE
        assign        iqPldWrPacket[2] = fab_chip.any.fabScalar.issueq.payloadRAM.data2wr_i;
      `endif
      `ifdef DISPATCH_FOUR_WIDE
        assign        iqPldWrPacket[3] = fab_chip.any.fabScalar.issueq.payloadRAM.data3wr_i;
      `endif
      `ifdef DISPATCH_FIVE_WIDE
        assign        iqPldWrPacket[4] = fab_chip.any.fabScalar.issueq.payloadRAM.data4wr_i;
      `endif
      `ifdef DISPATCH_SIX_WIDE
        assign        iqPldWrPacket[5] = fab_chip.any.fabScalar.issueq.payloadRAM.data5wr_i;
      `endif
      `ifdef DISPATCH_SEVEN_WIDE
        assign        iqPldWrPacket[6] = fab_chip.any.fabScalar.issueq.payloadRAM.data6wr_i;
      `endif
      `ifdef DISPATCH_EIGHT_WIDE
        assign        iqPldWrPacket[7] = fab_chip.any.fabScalar.issueq.payloadRAM.data7wr_i;
      `endif
      
      
      payloadPkt                                    iqPldRdPacket [0:`ISSUE_WIDTH-1];
        assign        iqPldRdPacket[0] = fab_chip.any.fabScalar.issueq.payloadRAM.data0_o;
      `ifdef ISSUE_TWO_WIDE
        assign        iqPldRdPacket[1] = fab_chip.any.fabScalar.issueq.payloadRAM.data1_o;
      `endif
      `ifdef ISSUE_THREE_WIDE
        assign        iqPldRdPacket[2] = fab_chip.any.fabScalar.issueq.payloadRAM.data2_o;
      `endif
      `ifdef ISSUE_FOUR_WIDE
        assign        iqPldRdPacket[3] = fab_chip.any.fabScalar.issueq.payloadRAM.data3_o;
      `endif
      `ifdef ISSUE_FIVE_WIDE
        assign        iqPldRdPacket[4] = fab_chip.any.fabScalar.issueq.payloadRAM.data4_o;
      `endif
      `ifdef ISSUE_SIX_WIDE
        assign        iqPldRdPacket[5] = fab_chip.any.fabScalar.issueq.payloadRAM.data5_o;
      `endif
      `ifdef ISSUE_SEVEN_WIDE
        assign        iqPldRdPacket[6] = fab_chip.any.fabScalar.issueq.payloadRAM.data6_o;
      `endif
      `ifdef ISSUE_EIGHT_WIDE
        assign        iqPldRdPacket[7] = fab_chip.any.fabScalar.issueq.payloadRAM.data7_o;
      `endif
      
      
      payloadPkt  [0:`ISSUE_WIDTH-1]                    rrPacket_l1;
      bypassPkt   [0:`ISSUE_WIDTH-1]                    bypassPacket;
      
      assign        rrPacket_l1                 = fab_chip.any.fabScalar.iq_regread.rrPacket_o;
      assign        bypassPacket                = fab_chip.any.fabScalar.registerfile.bypassPacket_i;
      
      fuPkt                           exePacket      [0:`ISSUE_WIDTH-1];
      fuPkt                           exePacket_s    [0:`ISSUE_WIDTH-1];
      fuPkt                           exePacket_c    [0:`ISSUE_WIDTH-1];
      
      
      assign    exePacket[0]      = fab_chip.any.fabScalar.exePipe0.execute.exePacket_i;
      assign    exePacket[1]      = fab_chip.any.fabScalar.exePipe1.execute.exePacket_i;
      assign    exePacket[2]      = fab_chip.any.fabScalar.exePipe2.execute.exePacket_i;
      //assign    exePacket_s[2]    = fab_chip.any.fabScalar.exePipe2.execute.simple_complex.salu.exePacket_i;
      //assign    exePacket_c[2]    = fab_chip.any.fabScalar.exePipe2.execute.simple_complex.calu.exePacket_i;
      
      `ifdef ISSUE_FOUR_WIDE
      assign    exePacket[3]      = fab_chip.any.fabScalar.exePipe3.execute.exePacket_i;
      //assign    exePacket_s[3]    = fab_chip.any.fabScalar.exePipe2.execute.simple_complex.salu.exePacket_i;
      //assign    exePacket_c[3]    = fab_chip.any.fabScalar.exePipe2.execute.simple_complex.calu.exePacket_i;
      `endif
      `ifdef ISSUE_FIVE_WIDE
      assign    exePacket[4]      = fab_chip.any.fabScalar.exePipe4.execute.exePacket_i;
      `endif
      `ifdef ISSUE_SIX_WIDE
      assign    exePacket[5]      = fab_chip.any.fabScalar.exePipe5.execute.exePacket_i;
      `endif
      
      
      memPkt                         memPacket;
      
      wbPkt                          lsuWbPacket;
      ldVioPkt                       ldVioPacket;
      
      assign    memPacket         = fab_chip.any.fabScalar.exePipe0.memPacket_o;
      assign    lsuWbPacket       = fab_chip.any.fabScalar.lsu.wbPacket_o;
      assign    ldVioPacket       = fab_chip.any.fabScalar.lsu.ldVioPacket_o;
      
      ctrlPkt     [0:`ISSUE_WIDTH-1]                     ctrlPacket;
      commitPkt   [0:`COMMIT_WIDTH-1]                    amtPacket;
      
      assign       ctrlPacket     = fab_chip.any.fabScalar.activeList.ctrlPacket_i;
      assign       amtPacket      = fab_chip.any.fabScalar.activeList.amtPacket_o;
      
      
      
      alPkt                               dataAl          [0:`COMMIT_WIDTH-1];
      wire [`EXECUTION_FLAGS-1:0]         ctrlAl          [0:`COMMIT_WIDTH-1];
      wire [`COMMIT_WIDTH-1:0]            commitReady;
      wire                                violateBit  [0:`COMMIT_WIDTH-1];
      reg  [`SIZE_ACTIVELIST_LOG-1:0]     headAddr [0:`COMMIT_WIDTH-1];
      reg  [`SIZE_ACTIVELIST_LOG-1:0]     tailAddr [0:`COMMIT_WIDTH-1];
      
      assign dataAl[0] = fab_chip.any.fabScalar.activeList.activeList.data0_o;
      assign ctrlAl[0] = fab_chip.any.fabScalar.activeList.ctrlActiveList.data0_o;
      assign commitReady[0] = fab_chip.any.fabScalar.activeList.executedActiveList.data0_o;
      assign violateBit[0] = fab_chip.any.fabScalar.activeList.ldViolateVector.data0_o;
      assign headAddr[0] = fab_chip.any.fabScalar.activeList.activeList.addr0_i;
      assign tailAddr[0] = fab_chip.any.fabScalar.activeList.activeList.addr0wr_i;
      
      `ifdef COMMIT_TWO_WIDE
      assign dataAl[1] = fab_chip.any.fabScalar.activeList.activeList.data1_o;
      assign ctrlAl[1] = fab_chip.any.fabScalar.activeList.ctrlActiveList.data1_o;
      assign commitReady[1] = fab_chip.any.fabScalar.activeList.executedActiveList.data1_o;
      assign violateBit[1] = fab_chip.any.fabScalar.activeList.ldViolateVector.data1_o;
      assign headAddr[1] = fab_chip.any.fabScalar.activeList.activeList.addr1_i;
      assign tailAddr[1] = fab_chip.any.fabScalar.activeList.activeList.addr1wr_i;
      `endif
      
      `ifdef COMMIT_THREE_WIDE
      assign dataAl[2] = fab_chip.any.fabScalar.activeList.activeList.data2_o;
      assign ctrlAl[2] = fab_chip.any.fabScalar.activeList.ctrlActiveList.data2_o;
      assign commitReady[2] = fab_chip.any.fabScalar.activeList.executedActiveList.data2_o;
      assign violateBit[2] = fab_chip.any.fabScalar.activeList.ldViolateVector.data2_o;
      assign headAddr[2] = fab_chip.any.fabScalar.activeList.activeList.addr2_i;
      assign tailAddr[2] = fab_chip.any.fabScalar.activeList.activeList.addr2wr_i;
      `endif
      
      `ifdef COMMIT_FOUR_WIDE
      assign dataAl[3] = fab_chip.any.fabScalar.activeList.activeList.data3_o;
      assign ctrlAl[3] = fab_chip.any.fabScalar.activeList.ctrlActiveList.data3_o;
      assign commitReady[3] = fab_chip.any.fabScalar.activeList.executedActiveList.data3_o;
      assign violateBit[3] = fab_chip.any.fabScalar.activeList.ldViolateVector.data3_o;
      assign headAddr[3] = fab_chip.any.fabScalar.activeList.activeList.addr3_i;
      assign tailAddr[3] = fab_chip.any.fabScalar.activeList.activeList.addr3wr_i;
      `endif
      
      reg                                 violateFlag [0:`COMMIT_WIDTH-1];
      reg                                 mispredFlag [0:`COMMIT_WIDTH-1];
      reg                                 exceptionFlag  [0:`COMMIT_WIDTH-1];
      
      always_comb
      begin
      	int i;
      	for (i = 0; i < `COMMIT_WIDTH; i = i + 1)
      	begin
      	/* The violate flag is used to mark a load violation.
      	 * An instruction with the violate bit set waits until it reaches 
      	 * the head of the AL and then causes a recovery without committing. */
      		violateFlag[i]    = violateBit[i] && commitReady[i];
      
      	/* The mispredict flag is used to mark a misprediction.
      	 * An instruction with the mispredict bit set commits only at 
      	 * the head of the AL. */
      		mispredFlag[i]    = ctrlAl[i][0] && commitReady[i];
      
      	/* The exception flag is used to mark the system call. 
      	 * An instruction with the exception bit set waits until it reaches 
      	 * the head of the AL before committing. After it has committed, 
      	 * a recovery occurs and the system call is handled. */
      		exceptionFlag[i]  = ctrlAl[i][1] && commitReady[i];
      	end
      	violateFlag[0]    = (violateBit[0] && commitReady[0]) || 
              (violateBit[1] && commitReady[0] && commitReady[1] && ctrlAl[0][3]);
      end
      
      
      always_ff @(posedge clk)
      begin : UPDATE_PHYSICAL_REG
          int i;
          for (i = 0; i < `ISSUE_WIDTH; i++)
          begin
              if (bypassPacket[i].valid)
              begin
                  PHYSICAL_REG[bypassPacket[i].tag] <= bypassPacket[i].data;
              end
          end
      end
      
      integer skip_instructions = 69;
      always_comb
      begin:COMMIT
      	int i;
      	reg [`COMMIT_WIDTH-1:0]        commitVector_f;
        reg [`COMMIT_WIDTH-1:0]        commitFission;
        reg [`SIZE_ACTIVELIST_LOG:0]   alCount;
        reg [`COMMIT_WIDTH-1:0]        commitVector;
        reg [`COMMIT_WIDTH-1:0]        commitVector_t1;
      
        alCount = fab_chip.any.fabScalar.activeList.activeListCnt_o;
      
      	totalCommit          = 0;
      
      	for (i = 0; i < `COMMIT_WIDTH; i = i + 1) 
      	begin
      		commitFission[i]  = ctrlAl[i][3] && commitReady[i];
      	end
      
      
      	commitVector_f[0] = (alCount > 0) & commitReady[0] & ~violateFlag[0]    & ~exceptionFlag[0];
      
      	for (i = 1; i < `COMMIT_WIDTH; i = i + 1) 
      	begin
      		commitVector_f[i] = (alCount > i) & commitReady[i] & ~mispredFlag[i] & ~mispredFlag[0] &
      		                     ~violateFlag[i] & ~exceptionFlag[i];
      	end
      
      	/* Retire the fission instructions together */
      	for (i = 0; i < `COMMIT_WIDTH-1; i = i + 1) 
      	begin
      		if (commitFission[i])
      		begin
      			commitVector[i] = commitVector_f[i] & commitVector_f[i+1] ;
      		end
      		else
      		begin
      			commitVector[i] = commitVector_f[i];
      		end
      	end
      
      	if (commitFission[`COMMIT_WIDTH-1])
      	begin
      		commitVector[`COMMIT_WIDTH-1] = 1'b0;
      	end
      	else
      	begin
      		commitVector[`COMMIT_WIDTH-1] = commitVector_f[`COMMIT_WIDTH-1];
      	end
      
      
        // Although the COMMIT_READY ram read port for a particular
        // RAM is already gated and the ready bit will 0 for an inactive
        // lane, it is better to put this mask here in case the RAMs are
        // power gated and logic levels are not guaranteed.
      `ifdef DYNAMIC_CONFIG
        commitVector = commitVector & commitLaneActive;
      `endif
      
      	commitVector_t1               = 4'h0;
      
        // May 19th - Rewritten the logic to make it per lane
        // RBRC
        // Extending to 4 bits
        casez ({{4-`COMMIT_WIDTH{1'b0}},commitVector})
          4'b0000:  begin
          end
          4'b??01:  begin
            commitVector_t1 = 4'h1;
            totalCommit     = 1;
          end
      `ifdef COMMIT_TWO_WIDE
          4'b?011:  begin
            commitVector_t1 = 4'h3;
            totalCommit     = 2;
          end
      `endif    
      `ifdef COMMIT_THREE_WIDE
          4'b0111:  begin
            commitVector_t1 = 4'h7;
            totalCommit     = 3;
          end
      `endif    
      `ifdef COMMIT_FOUR_WIDE
          4'b1111:  begin
            commitVector_t1 = 4'hf;
            totalCommit     = 4;
          end
      `endif    
          default: begin
            commitVector_t1 = 4'h0;
            totalCommit     = 0;
          end
        endcase
      end




`else //PNR_SIM



      logic [`ICACHE_LINE_SIZE-1:0][`ICACHE_NUM_LINES-1:0]                        data_array;
      logic [(`ICACHE_TAG_BITS*`ICACHE_INSTS_IN_LINE)-1:0][`ICACHE_NUM_LINES-1:0] tag_array;
  
      //assign  data_array = fab_chip.fabScalar.fs1.l1icache.icache.data_array; 
      //assign  tag_array  = fab_chip.fabScalar.fs1.l1icache.icache.tag_array; 

      fs2Pkt  [0:`FETCH_WIDTH-1]                   fs2Packet;
      fs2Pkt  [0:`FETCH_WIDTH-1]                   fs2Packet_l1;
      
      assign        fs2Packet     = fab_chip.fabScalar.fs1fs2.fs2Packet_i;
      assign        fs2Packet_l1  = fab_chip.fabScalar.fs1fs2.fs2Packet_o;
      
      decPkt  [0:`FETCH_WIDTH-1]                   decPacket;
      decPkt  [0:`FETCH_WIDTH-1]                   decPacket_l1;
      renPkt  [0:2*`FETCH_WIDTH-1]                 ibPacket;
      
      assign        decPacket     = fab_chip.fabScalar.fs2dec.decPacket_i;
      assign        decPacket_l1  = fab_chip.fabScalar.fs2dec.decPacket_o;
      assign        ibPacket      = fab_chip.fabScalar.decode.ibPacket_o;
      
      renPkt  [0:`DISPATCH_WIDTH-1]                renPacket;
      renPkt  [0:`DISPATCH_WIDTH-1]                renPacket_l1;
      
      assign        renPacket     = fab_chip.fabScalar.instBufRen.renPacket_i;
      assign        renPacket_l1  = fab_chip.fabScalar.instBufRen.renPacket_o;
      
      
      disPkt  [0:`DISPATCH_WIDTH-1]                     disPacket_l1;
      iqPkt   [0:`DISPATCH_WIDTH-1]                     iqPacket;
      alPkt   [0:`DISPATCH_WIDTH-1]                     alPacket;
      lsqPkt  [0:`DISPATCH_WIDTH-1]                     lsqPacket;
      
      assign        disPacket_l1                = fab_chip.fabScalar.renDis.disPacket_o;
      assign        iqPacket                    = fab_chip.fabScalar.dispatch.iqPacket_o;
      assign        alPacket                    = fab_chip.fabScalar.dispatch.alPacket_o;
      assign        lsqPacket                   = fab_chip.fabScalar.lsu.lsqPacket_i;
      
      iqEntryPkt    [0:`ISSUE_WIDTH-1]              iqGrantedEntry;
      iqEntryPkt    [0:`ISSUE_WIDTH-1]              iqFreedEntry  ;
      iqEntryPkt    [0:`DISPATCH_WIDTH-1]           iqFreeEntry   ;
      
      assign        iqGrantedEntry                = fab_chip.fabScalar.issueq.issueQfreelist.grantedEntry_i;
      assign        iqFreedEntry                  = fab_chip.fabScalar.issueq.issueQfreelist.freedEntry_o;
      assign        iqFreeEntry                   = fab_chip.fabScalar.issueq.issueQfreelist.freeEntry_o;
      
      payloadPkt                                    iqPldWrPacket [0:`DISPATCH_WIDTH-1];
        assign        iqPldWrPacket[0] = fab_chip.fabScalar.issueq.payloadRAM.data0wr_i;
      `ifdef DISPATCH_TWO_WIDE
        assign        iqPldWrPacket[1] = fab_chip.fabScalar.issueq.payloadRAM.data1wr_i;
      `endif
      `ifdef DISPATCH_THREE_WIDE
        assign        iqPldWrPacket[2] = fab_chip.fabScalar.issueq.payloadRAM.data2wr_i;
      `endif
      `ifdef DISPATCH_FOUR_WIDE
        assign        iqPldWrPacket[3] = fab_chip.fabScalar.issueq.payloadRAM.data3wr_i;
      `endif
      `ifdef DISPATCH_FIVE_WIDE
        assign        iqPldWrPacket[4] = fab_chip.fabScalar.issueq.payloadRAM.data4wr_i;
      `endif
      `ifdef DISPATCH_SIX_WIDE
        assign        iqPldWrPacket[5] = fab_chip.fabScalar.issueq.payloadRAM.data5wr_i;
      `endif
      `ifdef DISPATCH_SEVEN_WIDE
        assign        iqPldWrPacket[6] = fab_chip.fabScalar.issueq.payloadRAM.data6wr_i;
      `endif
      `ifdef DISPATCH_EIGHT_WIDE
        assign        iqPldWrPacket[7] = fab_chip.fabScalar.issueq.payloadRAM.data7wr_i;
      `endif
      
      
      payloadPkt                                    iqPldRdPacket [0:`ISSUE_WIDTH-1];
        assign        iqPldRdPacket[0] = fab_chip.fabScalar.issueq.payloadRAM.data0_o;
      `ifdef ISSUE_TWO_WIDE
        assign        iqPldRdPacket[1] = fab_chip.fabScalar.issueq.payloadRAM.data1_o;
      `endif
      `ifdef ISSUE_THREE_WIDE
        assign        iqPldRdPacket[2] = fab_chip.fabScalar.issueq.payloadRAM.data2_o;
      `endif
      `ifdef ISSUE_FOUR_WIDE
        assign        iqPldRdPacket[3] = fab_chip.fabScalar.issueq.payloadRAM.data3_o;
      `endif
      `ifdef ISSUE_FIVE_WIDE
        assign        iqPldRdPacket[4] = fab_chip.fabScalar.issueq.payloadRAM.data4_o;
      `endif
      `ifdef ISSUE_SIX_WIDE
        assign        iqPldRdPacket[5] = fab_chip.fabScalar.issueq.payloadRAM.data5_o;
      `endif
      `ifdef ISSUE_SEVEN_WIDE
        assign        iqPldRdPacket[6] = fab_chip.fabScalar.issueq.payloadRAM.data6_o;
      `endif
      `ifdef ISSUE_EIGHT_WIDE
        assign        iqPldRdPacket[7] = fab_chip.fabScalar.issueq.payloadRAM.data7_o;
      `endif
      
      
      payloadPkt  [0:`ISSUE_WIDTH-1]                    rrPacket_l1;
      bypassPkt   [0:`ISSUE_WIDTH-1]                    bypassPacket;
      
      assign        rrPacket_l1                 = fab_chip.fabScalar.iq_regread.rrPacket_o;
      assign        bypassPacket                = fab_chip.fabScalar.registerfile.bypassPacket_i;
      
      fuPkt                           exePacket      [0:`ISSUE_WIDTH-1];
      fuPkt                           exePacket_s    [0:`ISSUE_WIDTH-1];
      fuPkt                           exePacket_c    [0:`ISSUE_WIDTH-1];
      
      
      assign    exePacket[0]      = fab_chip.fabScalar.exePipe0.execute.exePacket_i;
      assign    exePacket[1]      = fab_chip.fabScalar.exePipe1.execute.exePacket_i;
      assign    exePacket[2]      = fab_chip.fabScalar.exePipe2.execute.exePacket_i;
      assign    exePacket_s[2]    = fab_chip.fabScalar.exePipe2.execute.simple_complex_salu.exePacket_i;
      assign    exePacket_c[2]    = fab_chip.fabScalar.exePipe2.execute.simple_complex_calu.exePacket_i;
      
      `ifdef ISSUE_FOUR_WIDE
      assign    exePacket[3]      = fab_chip.fabScalar.exePipe3.execute.exePacket_i;
      //assign    exePacket_s[3]    = fab_chip.fabScalar.exePipe2.execute.simple_complex_salu.exePacket_i;
      //assign    exePacket_c[3]    = fab_chip.fabScalar.exePipe2.execute.simple_complex_calu.exePacket_i;
      `endif
      `ifdef ISSUE_FIVE_WIDE
      assign    exePacket[4]      = fab_chip.fabScalar.exePipe4.execute.exePacket_i;
      `endif
      `ifdef ISSUE_SIX_WIDE
      assign    exePacket[5]      = fab_chip.fabScalar.exePipe5.execute.exePacket_i;
      `endif
      
      
      memPkt                         memPacket;
      
      wbPkt                          lsuWbPacket;
      ldVioPkt                       ldVioPacket;
      
      assign    memPacket         = fab_chip.fabScalar.exePipe0.memPacket_o;
      assign    lsuWbPacket       = fab_chip.fabScalar.lsu.wbPacket_o;
      assign    ldVioPacket       = fab_chip.fabScalar.lsu.ldVioPacket_o;
      
      ctrlPkt     [0:`ISSUE_WIDTH-1]                     ctrlPacket;
      commitPkt   [0:`COMMIT_WIDTH-1]                    amtPacket;
      
      assign       ctrlPacket     = fab_chip.fabScalar.activeList.ctrlPacket_i;
      assign       amtPacket      = fab_chip.fabScalar.activeList.amtPacket_o;
      
      
      
      alPkt                               dataAl          [0:`COMMIT_WIDTH-1];
      wire [`EXECUTION_FLAGS-1:0]         ctrlAl          [0:`COMMIT_WIDTH-1];
      wire [`COMMIT_WIDTH-1:0]            commitReady;
      wire                                violateBit  [0:`COMMIT_WIDTH-1];
      reg  [`SIZE_ACTIVELIST_LOG-1:0]     headAddr [0:`COMMIT_WIDTH-1];
      reg  [`SIZE_ACTIVELIST_LOG-1:0]     tailAddr [0:`COMMIT_WIDTH-1];
      
      assign dataAl[0] = fab_chip.fabScalar.activeList.activeList.data0_o;
      assign ctrlAl[0] = fab_chip.fabScalar.activeList.ctrlActiveList.data0_o;
      assign commitReady[0] = fab_chip.fabScalar.activeList.executedActiveList.data0_o;
      assign violateBit[0] = fab_chip.fabScalar.activeList.ldViolateVector.data0_o;
      assign headAddr[0] = fab_chip.fabScalar.activeList.activeList.addr0_i;
      assign tailAddr[0] = fab_chip.fabScalar.activeList.activeList.addr0wr_i;
      
      `ifdef COMMIT_TWO_WIDE
      assign dataAl[1] = fab_chip.fabScalar.activeList.activeList.data1_o;
      assign ctrlAl[1] = fab_chip.fabScalar.activeList.ctrlActiveList.data1_o;
      assign commitReady[1] = fab_chip.fabScalar.activeList.executedActiveList.data1_o;
      assign violateBit[1] = fab_chip.fabScalar.activeList.ldViolateVector.data1_o;
      assign headAddr[1] = fab_chip.fabScalar.activeList.activeList.addr1_i;
      assign tailAddr[1] = fab_chip.fabScalar.activeList.activeList.addr1wr_i;
      `endif
      
      `ifdef COMMIT_THREE_WIDE
      assign dataAl[2] = fab_chip.fabScalar.activeList.activeList.data2_o;
      assign ctrlAl[2] = fab_chip.fabScalar.activeList.ctrlActiveList.data2_o;
      assign commitReady[2] = fab_chip.fabScalar.activeList.executedActiveList.data2_o;
      assign violateBit[2] = fab_chip.fabScalar.activeList.ldViolateVector.data2_o;
      assign headAddr[2] = fab_chip.fabScalar.activeList.activeList.addr2_i;
      assign tailAddr[2] = fab_chip.fabScalar.activeList.activeList.addr2wr_i;
      `endif
      
      `ifdef COMMIT_FOUR_WIDE
      assign dataAl[3] = fab_chip.fabScalar.activeList.activeList.data3_o;
      assign ctrlAl[3] = fab_chip.fabScalar.activeList.ctrlActiveList.data3_o;
      assign commitReady[3] = fab_chip.fabScalar.activeList.executedActiveList.data3_o;
      assign violateBit[3] = fab_chip.fabScalar.activeList.ldViolateVector.data3_o;
      assign headAddr[3] = fab_chip.fabScalar.activeList.activeList.addr3_i;
      assign tailAddr[3] = fab_chip.fabScalar.activeList.activeList.addr3wr_i;
      `endif
      
      reg                                 violateFlag [0:`COMMIT_WIDTH-1];
      reg                                 mispredFlag [0:`COMMIT_WIDTH-1];
      reg                                 exceptionFlag  [0:`COMMIT_WIDTH-1];
      
      always_comb
      begin
      	int i;
      	for (i = 0; i < `COMMIT_WIDTH; i = i + 1)
      	begin
      	/* The violate flag is used to mark a load violation.
      	 * An instruction with the violate bit set waits until it reaches 
      	 * the head of the AL and then causes a recovery without committing. */
      		violateFlag[i]    = violateBit[i] && commitReady[i];
      
      	/* The mispredict flag is used to mark a misprediction.
      	 * An instruction with the mispredict bit set commits only at 
      	 * the head of the AL. */
      		mispredFlag[i]    = ctrlAl[i][0] && commitReady[i];
      
      	/* The exception flag is used to mark the system call. 
      	 * An instruction with the exception bit set waits until it reaches 
      	 * the head of the AL before committing. After it has committed, 
      	 * a recovery occurs and the system call is handled. */
      		exceptionFlag[i]  = ctrlAl[i][1] && commitReady[i];
      	end
      	violateFlag[0]    = (violateBit[0] && commitReady[0]) || 
              (violateBit[1] && commitReady[0] && commitReady[1] && ctrlAl[0][3]);
      end
      
      
      always_ff @(posedge clk)
      begin : UPDATE_PHYSICAL_REG
          int i;
          for (i = 0; i < `ISSUE_WIDTH; i++)
          begin
              if (bypassPacket[i].valid)
              begin
                  PHYSICAL_REG[bypassPacket[i].tag] <= bypassPacket[i].data;
              end
          end
      end
      
      integer skip_instructions = 69;
      always_comb
      begin:COMMIT
      	int i;
      	reg [`COMMIT_WIDTH-1:0]        commitVector_f;
        reg [`COMMIT_WIDTH-1:0]        commitFission;
        reg [`SIZE_ACTIVELIST_LOG:0]   alCount;
        reg [`COMMIT_WIDTH-1:0]        commitVector;
        reg [`COMMIT_WIDTH-1:0]        commitVector_t1;
      
        alCount = fab_chip.fabScalar.activeList.activeListCnt_o;
      
      	totalCommit          = 0;
      
      	for (i = 0; i < `COMMIT_WIDTH; i = i + 1) 
      	begin
      		commitFission[i]  = ctrlAl[i][3] && commitReady[i];
      	end
      
      
      	commitVector_f[0] = (alCount > 0) & commitReady[0] & ~violateFlag[0]    & ~exceptionFlag[0];
      
      	for (i = 1; i < `COMMIT_WIDTH; i = i + 1) 
      	begin
      		commitVector_f[i] = (alCount > i) & commitReady[i] & ~mispredFlag[i] & ~mispredFlag[0] &
      		                     ~violateFlag[i] & ~exceptionFlag[i];
      	end
      
      	/* Retire the fission instructions together */
      	for (i = 0; i < `COMMIT_WIDTH-1; i = i + 1) 
      	begin
      		if (commitFission[i])
      		begin
      			commitVector[i] = commitVector_f[i] & commitVector_f[i+1] ;
      		end
      		else
      		begin
      			commitVector[i] = commitVector_f[i];
      		end
      	end
      
      	if (commitFission[`COMMIT_WIDTH-1])
      	begin
      		commitVector[`COMMIT_WIDTH-1] = 1'b0;
      	end
      	else
      	begin
      		commitVector[`COMMIT_WIDTH-1] = commitVector_f[`COMMIT_WIDTH-1];
      	end
      
      
        // Although the COMMIT_READY ram read port for a particular
        // RAM is already gated and the ready bit will 0 for an inactive
        // lane, it is better to put this mask here in case the RAMs are
        // power gated and logic levels are not guaranteed.
      `ifdef DYNAMIC_CONFIG
        commitVector = commitVector & commitLaneActive;
      `endif
      
      	commitVector_t1               = 4'h0;
      
        // May 19th - Rewritten the logic to make it per lane
        // RBRC
        // Extending to 4 bits
        casez ({{4-`COMMIT_WIDTH{1'b0}},commitVector})
          4'b0000:  begin
          end
          4'b??01:  begin
            commitVector_t1 = 4'h1;
            totalCommit     = 1;
          end
      `ifdef COMMIT_TWO_WIDE
          4'b?011:  begin
            commitVector_t1 = 4'h3;
            totalCommit     = 2;
          end
      `endif    
      `ifdef COMMIT_THREE_WIDE
          4'b0111:  begin
            commitVector_t1 = 4'h7;
            totalCommit     = 3;
          end
      `endif    
      `ifdef COMMIT_FOUR_WIDE
          4'b1111:  begin
            commitVector_t1 = 4'hf;
            totalCommit     = 4;
          end
      `endif    
          default: begin
            commitVector_t1 = 4'h0;
            totalCommit     = 0;
          end
        endcase
      end

`endif //PNR_SIM


//`ifdef VERIFY_COMMIT
always @(posedge clk)
begin: VERIFY_INSTRUCTIONS
    reg [`SIZE_PC-1:0]           PC           [`COMMIT_WIDTH-1:0];
    reg [`SIZE_RMT_LOG-1:0]      logDest      [`COMMIT_WIDTH-1:0];
    reg [`SIZE_PHYSICAL_LOG-1:0] phyDest      [`COMMIT_WIDTH-1:0];
    reg [`SIZE_DATA-1:0]         result       [`COMMIT_WIDTH-1:0];
    reg                          isBranch     [`COMMIT_WIDTH-1:0];
    reg                          isMispredict [`COMMIT_WIDTH-1:0];
    reg                          eChecker     [`COMMIT_WIDTH-1:0];
    reg                          isFission    [`COMMIT_WIDTH-1:0];
    reg [`SIZE_PC-1:0]           lastCommitPC;
    int i;


    for (i = 0; i < `COMMIT_WIDTH; i++)
    begin
        PC[i]           = dataAl[i].pc;
        logDest[i]      = dataAl[i].logDest;
        phyDest[i]      = dataAl[i].phyDest;
        result[i]       = PHYSICAL_REG[phyDest[i]];
  
        eChecker[i]     = (totalCommit >= (i+1)) ? 1'h1 : 1'h0;
        isFission[i]    = ctrlAl[i][3] & commitReady[i];
        isBranch[i]     = ctrlAl[i][5];

        isMispredict[i] = ctrlAl[i][0] & ctrlAl[i][5];
    end

    if (eChecker[0] && (skip_instructions != 0) && verifyCommits)
    begin
        skip_instructions = skip_instructions - totalCommit;
    end

    else if(verifyCommits)
    begin
        if (lastCommitPC == PC[0] && eChecker[0])
        begin
            lastCommitPC = PC[0];
        end

        else
        begin
            if (eChecker[0]) lastCommitPC = PC[0];

            $getRetireInstPCNetSim(eChecker[0],CYCLE_COUNT,PC[0],logDest[0],result[0],isFission[0],0);
        end

    `ifdef COMMIT_TWO_WIDE
        if (lastCommitPC == PC[1] && eChecker[1])
        begin
            lastCommitPC = PC[1];
        end

        else
        begin
            if(eChecker[1]) lastCommitPC = PC[1];

            $getRetireInstPCNetSim(eChecker[1],CYCLE_COUNT,PC[1],logDest[1],result[1],isFission[1],1);
        end
    `endif

    `ifdef COMMIT_THREE_WIDE
        if (lastCommitPC == PC[2] && eChecker[2])
        begin
            lastCommitPC = PC[2];
        end

        else
        begin
            if(eChecker[2]) lastCommitPC = PC[2];

            $getRetireInstPCNetSim(eChecker[2],CYCLE_COUNT,PC[2],logDest[2],result[2],isFission[2],1);
        end
    `endif

    `ifdef COMMIT_FOUR_WIDE
        if (lastCommitPC == PC[3] && eChecker[3])
        begin
            lastCommitPC = PC[3];
        end

        else
        begin
            if(eChecker[3]) lastCommitPC = PC[3];

            $getRetireInstPCNetSim(eChecker[3],CYCLE_COUNT,PC[3],logDest[3],result[3],isFission[3],1);
        end
    `endif
    end
end
//`endif

task copyRF;

    integer i;

    begin
        for (i = 0; i < 34; i++)
        begin
            //fabScalar.registerfile.PhyRegFile_byte0.ram[i] = LOGICAL_REG[i][7:0];
            //fabScalar.registerfile.PhyRegFile_byte1.ram[i] = LOGICAL_REG[i][15:8];
            //fabScalar.registerfile.PhyRegFile_byte2.ram[i] = LOGICAL_REG[i][23:16];
            //fabScalar.registerfile.PhyRegFile_byte3.ram[i] = LOGICAL_REG[i][31:24];
        end

    end
endtask

task copySimRF;

    int i;

    begin
        for (i = 0; i < 34; i++)
        begin
            PHYSICAL_REG[i] = LOGICAL_REG[i];
        end

        for (i = 34; i < `SIZE_PHYSICAL_TABLE; i++)
        begin
            PHYSICAL_REG[i] = 0;
        end
    end
endtask

task init_registers;
    integer i;
    reg  [31:0] opcode;
    reg  [7:0]  dest;
    reg  [7:0]  src1;
    reg  [7:0]  src2;
    reg  [15:0] immed;
    reg  [25:0] target; 

    begin
        for (i = 1; i < 34; i = i + 1)
        begin
            opcode  = {24'h0, `LUI};
            dest    = i;
            immed   = LOGICAL_REG[i][31:16];
            `WRITE_WORD(opcode, (32'h0000_0000 + 16*(i-1)));
            `WRITE_WORD({8'h0, dest, immed}, (32'h0000_0000 + 16*(i-1)+4));
            $display("LUI = Opcode: %x dest: %x immed: %x addr: %x",opcode,dest,immed,(32'h0000_0000 + 16*(i-1)));

            opcode  = {24'h0, `ORI};
            dest    = i;
            src1    = i;
            immed   = LOGICAL_REG[i][15:0];
            `WRITE_WORD(opcode, (32'h0000_0000 + 16*(i-1)+8)); 
            `WRITE_WORD({src1, dest, immed}, (32'h0000_0000 + 16*(i-1)+12)); 
            /* $display("@%d[%08x]", i, LOGICAL_REG[i]); */
            PHYSICAL_REG[i] = LOGICAL_REG[i];
            $display("ORI = Opcode: %x dest: %x src1: %x immed: %x addr: %x",opcode,dest,src1,immed,(32'h0000_0000 + 16*(i-1)+2));
        end

        // return from subroutine
        opcode  = {24'h0, `RET};
        target  = `GET_ARCH_PC >> 2;
        `WRITE_WORD(opcode, (32'h0000_0000 + 16*(i-1))); 
        `WRITE_WORD({6'h0, target}, (32'h0000_0000 + 16*(i-1)+4)); 

        // skip two instructions per register plus 1 for jump
        skip_instructions = 2*33 + 1;
    end
endtask

task load_kernel_scratch;
 integer  ram_index;
 integer  offset;
 integer  data_file; 
 integer  scan_file; 

  $display("Loading ICACHE data\n");
  for(ram_index = 0; ram_index < (2**(`ICACHE_INDEX_BITS+`ICACHE_BYTES_IN_LINE_LOG)) ; ram_index++)
  begin
    //instScratchAddr   = {offset[2:0],ram_index[7:0]};
    #(IO_CLKPERIOD);
    regAddr   = 6'h30;
    regWrData = ram_index[7:0]; 
    regWrEn   = 1'b1;
    #(IO_CLKPERIOD);
    regAddr   = 6'h31;
    regWrData = ram_index[`ICACHE_INDEX_BITS+`ICACHE_BYTES_IN_LINE_LOG-1:8]; 
    regWrEn   = 1'b1;
    #(IO_CLKPERIOD);
    regAddr   = 6'h32;
    regWrData = ram_index[7:0]-2;
    regWrEn   = 1'b1;
//      regWrData = kernel_line[8*(offset+1)-1-:8];
    #(IO_CLKPERIOD);
    regWrEn   = 1'b0;
  end

endtask
  
task read_kernel_scratch;
 integer  ram_index;
 integer  offset;
 integer  data_file; 
 integer  scan_file; 
 reg  [7:0] check_data;

  $display("Reading ICACHE data\n");
  for(ram_index = 0; ram_index < (2**(`ICACHE_INDEX_BITS+`ICACHE_BYTES_IN_LINE_LOG)) ; ram_index++)
  begin
    regAddr   = 6'h30;    // Address LSB
    regWrData = ram_index[7:0]; 
    regWrEn   = 1'b1;
    #(IO_CLKPERIOD);
    regAddr   = 6'h31;    // Address MSB
    regWrData = ram_index[`ICACHE_INDEX_BITS+`ICACHE_BYTES_IN_LINE_LOG-1:8]; 
    regWrEn   = 1'b1;
    #(IO_CLKPERIOD);
    regWrEn   = 1'b0;
    #(3*IO_CLKPERIOD);  // Takes 2 cycles for data to be read and synchronized
    regAddr   = 6'h33;  // Issue indirect read address
    #(IO_CLKPERIOD);
    check_data = ram_index[7:0] - 2'h2;
    if(regRdData != check_data)
    begin
      $display("Cycle: %0d ICACHE READ MISMATCH at index %03x \n",CYCLE_COUNT,ram_index);
      $display("Read %02x , expected %02x\n",regRdData,(ram_index[7:0] - 2));
    end
  end
endtask

task load_data_scratch;
 integer  ram_index;
 integer  offset;
 integer  data_file; 
 integer  scan_file; 

  $display("Loading DCACHE data\n");
  for(ram_index = 0; ram_index < (2**(`DCACHE_INDEX_BITS+`DCACHE_BYTES_IN_LINE_LOG)) ; ram_index++)
  begin
    //instScratchAddr   = {offset[2:0],ram_index[7:0]};
    #(IO_CLKPERIOD);
    regAddr   = 6'h34;
    regWrData = ram_index[7:0]; 
    regWrEn   = 1'b1;
    #(IO_CLKPERIOD);
    regAddr   = 6'h35;
    regWrData = ram_index[`DCACHE_INDEX_BITS+`DCACHE_BYTES_IN_LINE_LOG-1:8]; 
    regWrEn   = 1'b1;
    #(IO_CLKPERIOD);
    regAddr   = 6'h36;
    regWrData = ram_index[7:0]-2;
    regWrEn   = 1'b1;
//      regWrData = kernel_line[8*(offset+1)-1-:8];
    #(IO_CLKPERIOD);
    regWrEn   = 1'b0;
  end

endtask
  
task read_data_scratch;
 integer  ram_index;
 integer  offset;
 integer  data_file; 
 integer  scan_file; 
 reg  [`REG_DATA_WIDTH-1:0] check_data;

  $display("Reading DCACHE data\n");
  for(ram_index = 0; ram_index < (2**(`DCACHE_INDEX_BITS+`DCACHE_BYTES_IN_LINE_LOG)) ; ram_index++)
  begin
    regAddr   = 6'h34;    // Address LSB
    regWrData = ram_index[7:0]; 
    regWrEn   = 1'b1;
    #(IO_CLKPERIOD);
    regAddr   = 6'h35;    // Address MSB
    regWrData = ram_index[`DCACHE_INDEX_BITS+`DCACHE_BYTES_IN_LINE_LOG-1:8]; 
    regWrEn   = 1'b1;
    #(IO_CLKPERIOD);
    regWrEn   = 1'b0;
    #(3*IO_CLKPERIOD);  // Takes 2 cycles for data to be read and synchronized
    regAddr   = 6'h37;  // Issue indirect read address
    #(IO_CLKPERIOD);
    check_data = ram_index[7:0] - 2'h2;
    if(regRdData != check_data)
    begin
      $display("Cycle: %0d DCACHE READ MISMATCH at index %03x \n",CYCLE_COUNT,ram_index);
      $display("Read %02x , expected %02x\n",regRdData,(ram_index[7:0] - 2));
    end
  end
endtask

//task to load the PRF from checkpoint
task load_checkpoint_PRF;
  integer  ram_index;
  integer  offset;
  
  for(ram_index = 0; ram_index < `SIZE_PHYSICAL_TABLE ; ram_index++)
    begin
    for(offset = 0; offset < 4 ; offset++)
    begin
      debugPRFAddr      = {offset[`SIZE_DATA_BYTE_OFFSET-1:0],ram_index[`SIZE_PHYSICAL_LOG-1:0]};
      debugPRFWrEn      = 1;   
      debugPRFWrData    = offset+ram_index;
      #(2*CLKPERIOD);
    end
    end
  debugPRFWrEn      = 0;
endtask

//task to read the PRF byte by byte
task read_checkpoint_PRF;
  integer  ram_index;
  integer  offset;

  for(ram_index = 0; ram_index < `SIZE_PHYSICAL_TABLE ; ram_index++)
  begin
    for(offset = 3; offset >= 0 ; offset--)
    begin
      debugPRFAddr      = {offset[`SIZE_DATA_BYTE_OFFSET-1:0],ram_index[`SIZE_PHYSICAL_LOG-1:0]};
      //debugPRFWrEn      = 1;  
      #(2*CLKPERIOD);
      if(debugPRFRdData      != offset+ram_index)
      begin
        $display("READ MISMATCH at %x index %d byte\n",ram_index,offset);
        $display("Read %x , expected %x\n",debugPRFRdData,offset+ram_index);
      end
    end
  end
endtask

//task to read the ARF byte by byte
task read_PRF;
  integer  ram_index;
  integer  offset;
  reg  [7:0]      captureRF[3:0]; 

  for(ram_index = 0; ram_index < `SIZE_PHYSICAL_TABLE ; ram_index++)
    begin
    for(offset = 3; offset >= 0 ; offset--)
    begin
      regAddr   = 6'h30;    // Address LSB
      regWrData = {offset[`SIZE_DATA_BYTE_OFFSET-1:0],ram_index[`SIZE_PHYSICAL_LOG-1:0]}; 
      regWrEn   = 1'b1;
      #(2*IO_CLKPERIOD);
      captureRF[offset] = debugPRFRdData;
      if(offset == 0)
      $display("Phys Reg %02x read %x%x%x%x\n",ram_index,captureRF[3],captureRF[2],captureRF[1],captureRF[0]);
    end
  end
endtask

//task to read the ARF byte by byte
task read_AMT;
  integer  ram_index;

  for(ram_index = 0; ram_index < `SIZE_RMT ; ram_index++)
  begin
    regAddr   = 6'h38;   // Indirect Address Reg 
    regWrData = {{(8-`SIZE_RMT_LOG){1'b0}},ram_index[`SIZE_RMT_LOG-1:0]}; 
    regWrEn   = 1'b1;
    #(IO_CLKPERIOD);
    regWrEn   = 1'b0;
    #(IO_CLKPERIOD);
    regAddr   = 6'h39;   // Read AMT Data reg
    #(3*IO_CLKPERIOD);
    $display("Log Reg: %02x -> Phys Reg %2x\n", ram_index,regRdData);
  end
endtask


`ifdef SCRATCH_PAD

  task load_inst_scratch;
   integer  ram_index;
   integer  offset;
   
   for(ram_index = 0; ram_index < `DEBUG_INST_RAM_DEPTH ; ram_index++ )
   //for(ram_index = 0; ram_index < 2 ; ram_index++ )
    begin
    for(offset =0; offset < 5 ; offset ++)
    begin
      instScratchAddr   = {offset[2:0],ram_index[7:0]};
      instScratchWrEn   = 1;   
      instScratchWrData = ram_index[7:0]^offset[7:0];
      #(CLKPERIOD);
    end
    end
  endtask
  
  //task to load the INSTRUCTION scratch pad with the microbenchmark
//  task load_kernel_scratch;
//   integer  ram_index;
//   integer  offset;
//   integer  data_file; 
//   integer  scan_file; 
//   reg [`DEBUG_INST_RAM_WIDTH-1:0] kernel_line;
//  
//   data_file = $fopen("kernel.dat","r");
//  
//   for(ram_index = 0; ram_index < `DEBUG_INST_RAM_DEPTH ; ram_index++ )
//    begin
//    scan_file = $fscanf(data_file, "%10x\n",kernel_line);
//    for(offset = 0; offset < 5 ; offset ++)
//    begin
//      instScratchAddr   = {offset[2:0],ram_index[7:0]};
//      instScratchWrEn   = 1;   
//      instScratchWrData = kernel_line[8*(offset+1)-1-:8];
//      #(CLKPERIOD);
//    end
//    end
//  endtask
//  
  //task to read the INSTRUCTION scratch pad
  task read_inst_scratch;
   integer ram_index;
   integer offset;
  for(ram_index = 0; ram_index < `DEBUG_INST_RAM_DEPTH ; ram_index++ )
    begin
    for(offset =0; offset < 5 ; offset ++)
    begin
      instScratchAddr   = {offset[2:0],ram_index[7:0]};   
      #(CLKPERIOD);
      if(instScratchRdData != (ram_index[7:0]^offset[7:0]))
      begin
        $display("READ MISMATCH at %x index %d byte\n",ram_index,offset);
        $display("Read %x , expected %x\n",instScratchRdData,ram_index[7:0]^offset[7:0]);
      end
    end
   end
  endtask

  task load_data_scratch;
   integer  ram_index;
   integer  offset;
   integer  data_file; 
   integer  scan_file; 
   reg [`DEBUG_DATA_RAM_WIDTH-1:0] data_line;
  
   data_file = $fopen("data.dat","r");
  
   for(ram_index = 0; ram_index < `DEBUG_DATA_RAM_DEPTH ; ram_index++ )
    begin
    scan_file = $fscanf(data_file, "%8x\n",data_line);
    for(offset = 0; offset < 3 ; offset ++)
    begin
      dataScratchAddr   = {offset[1:0],ram_index[7:0]};
      dataScratchWrEn   = 1;   
      dataScratchWrData = data_line[8*(offset+1)-1-:8];
      #(CLKPERIOD);
    end
    end
  endtask
  
  task read_data_scratch;
   integer  ram_index;
   integer  offset;
   integer  data_file; 
   integer  scan_file; 
   reg [`DEBUG_DATA_RAM_WIDTH-1:0] data_line;
  
   data_file = $fopen("data.dat","r");
  for(ram_index = 0; ram_index < `DEBUG_DATA_RAM_DEPTH ; ram_index++ )
    begin
    scan_file = $fscanf(data_file, "%8x\n",data_line);
    for(offset =0; offset < 3 ; offset ++)
    begin
      dataScratchAddr   = {offset[1:0],ram_index[7:0]};   
      #(CLKPERIOD);
      //if(dataScratchRdData != data_line[8*(offset+1)-1-:8])
      if(dataScratchRdData != data_line[8*(offset+1)-1-:8])
      begin
        $display("READ MISMATCH at %x index %d byte\n",ram_index,offset);
        $display("Read %x , expected %x\n",dataScratchRdData,data_line[8*(offset+1)-1-:8]);
      end
    end
   end
  endtask
  
`endif // SCRATCH_PAD


  task scan_in_chain1;
   integer  scan_index;
   integer  dat_file; 
   integer  scan_file; 
   reg      scan_line;
   integer  scan_index_2;
   integer  dat_file_2; 
   integer  scan_file_2; 
   reg      scan_line_2;
  begin 
   dat_file = $fopen("scan_in.dat","r");
   dat_file_2 = $fopen("scan_in_2.dat","r");
  
   for(scan_index = 0; scan_index <= 11305; scan_index++ )
    begin
   	scan_file = $fscanf(dat_file, "%b", scan_line);
    scan_file_2 = $fscanf(dat_file_2, "%b", scan_line_2);
    	test_se  = 1'b1;   
	@( posedge data_source)
	begin
    	test_si1 = scan_line;
    	test_si2 = scan_line_2;
	end
   // 	data_source = 1'b0;
   // 	#(10);
   // 	data_source = 1'b1;
   // 	#(10);
    end
  end
  test_se  = 1'b0;   
 // scan_lookup();  
 // scan_lookup_2();  
  $display("I Did my job - Scan Chain 1\n");
  endtask

  task scan_out_chain1;
   integer  scan_index;
   integer  dat_file; 
   integer  scan_file; 
   reg      scan_line;
   integer  scan_index_2;
   integer  dat_file_2; 
   integer  scan_file_2; 
   reg      scan_line_2;
  begin
   dat_file = $fopen("scan_out.dat","w");
   dat_file_2 = $fopen("scan_out_2.dat","w");
   // scan_lookup();  
   // scan_lookup_2();  
    for(scan_index = 0; scan_index <= 11304; scan_index++ )
    begin
    	test_se  = 1'b1;   
	  @( posedge data_source)
	  begin
    	$fwrite(dat_file, "%b\n", test_so1);
    	$fwrite(dat_file_2, "%b\n", test_so2);
	  end
    //	data_source = 1'b1;
    //	#(10);
    //	data_source = 1'b0;
    //	#(10);
   end
  end
  test_se  = 1'b0;   
  $display("I Did my job - Scan Out\n");
  endtask
 
  task scan_in_chain2;
   integer  scan_index_2;
   integer  dat_file_2; 
   integer  scan_file_2; 
   reg      scan_line_2;
  begin 
   dat_file_2 = $fopen("scan_in_2.dat","r");
   for(scan_index_2 = 0; scan_index_2 <= 11304 ; scan_index_2++ )
    begin
    	scan_file_2 = $fscanf(dat_file_2, "%b", scan_line_2);
    //	scan_file = $fread(scan_line, dat_file);        
    //    $display("scan_index:%d scan_line:%b",scan_index, scan_line); 
    	test_se  = 1'b1;   
    	test_si2 = scan_line_2;
    	data_source = 1'b0;
    	#(10);
    	data_source = 1'b1;
    	#(10);
    end
  end
  test_se  = 1'b0;   
//  scan_lookup_2();  
  $display("I Did my job - Scan Chain 2\n");
  endtask

  task scan_out_chain2;
   integer  scan_index_2;
   integer  dat_file_2; 
   integer  scan_file_2; 
   reg      scan_line_2;
  begin
   dat_file_2 = $fopen("scan_out_2.dat","w");
 //  scan_lookup_2();  
    for(scan_index_2 = 0; scan_index_2 <= 11304 ; scan_index_2++ )
    begin
    	test_se  = 1'b1;   
    	$fwrite(dat_file_2, "%b\n", test_so2);
    	data_source = 1'b1;
    	#(10);
    	data_source = 1'b0;
    	#(10);
   end
  end
  endtask

`ifdef PERF_MON

task read_perf_mon;
  integer  index;
  
  //perfMonRegRun        = 1'b1;
  regWrEn   = 1'b1;
  regAddr   = 6'h1A;
  regWrData = 8'h01;  
  #CLKPERIOD;
  regWrEn   = 1'b0;
 
  #(1000*CLKPERIOD)

  //perfMonRegRun        = 1'b0;
  regWrEn   = 1'b1;
  regAddr   = 6'h1A;
  regWrData = 8'h00 ; 
  #CLKPERIOD;
  regWrEn   = 1'b0;

  for(index = 8'h00; index < 8'h05 ; index++ )
  begin
    //perfMonRegAddr       = index[7:0];
  regAddr   = 6'h19;
  regWrData = index[7:0] ;
  case(index)
  00:$display("Events : totalCycles   : "); 
  01:$display("Events : commitStore   : ");
  02:$display("Events : commitLoad    : ");
  03:$display("Events : recoverflag   : ");
  04:$display("Events : loadViolation   : "); 
  05:$display("Events : totalCommit     : ");
  endcase
  read_4_byte();
  end

  for(index = 8'h10; index < 8'h12 ; index++ )
  begin
  //  perfMonRegAddr       = index[7:0];
  regAddr   = 6'h19;
  regWrData = index[7:0] ; 
  case(index)
  8'h10:$display("Occupancy : ibCount,flCount,iqCount,ldqCount : ");
  8'h11:$display("Occupancy : LSB 16 bit -- stqCount,commitCount: ");
  endcase
  read_4_byte();
  end
  for(index = 8'h20; index < 8'h21 ; index++ )
  begin
  //  perfMonRegAddr       = index[7:0];
  regAddr   = 6'h19;
  regWrData = index[7:0] ;
  $display("LSB 9 bit -- program_status_word : "); 
  read_4_byte();
  end
  for(index = 8'h30; index < 8'h32 ; index++ )
  begin
  //  perfMonRegAddr       = index[7:0];
  regAddr   = 6'h19;
  regWrData = index[7:0] ; 
  case(index)
  8'h30:$display("fs1fs2Valid_count,fs2DecValid_count,renDisValid_count,instBufRenValid_countibCount : ");
  8'h31:$display("LSB 16 bit -- iqValid_count,iqRegReadValid_count  : ");
  endcase
  read_4_byte();
  end
  for(index = 8'h40; index < 8'h49 ; index++ )
  begin
  //  perfMonRegAddr       = index[7:0];
  regAddr   = 6'h19;
  regWrData = index[7:0] ;
  case(index)
  8'h40:$display("Events : fetch1_stall   : ");
  8'h41:$display("Events : ctiq_stall     : ");
  8'h42:$display("Events : instBuf_stall  : ");
  8'h43:$display("Events : freelist_stall : ");
  8'h44:$display("Events : backend_stall  : ");
  8'h45:$display("Events : ldq_stall      : ");
  8'h46:$display("Events : stq_stall      : ");
  8'h47:$display("Events : iq_stall       : ");
  8'h48:$display("Events : rob_stall      : ");     
  endcase 
  read_4_byte();
  end
  for(index = 8'h50; index < 8'h55 ; index++ )
  begin
  //  perfMonRegAddr       = index[7:0];
  regAddr   = 6'h19;
  regWrData = index[7:0] ;
  case(index)
  8'h50:$display("Events : instMiss   : ");
  8'h51:$display("Events : loadMiss     : ");
  8'h52:$display("Events : storeMiss  : ");
  8'h53:$display("Events : l2InstFetchReq : ");
  8'h54:$display("Events : l2DataFetchReq  : ");
  endcase 
  read_4_byte();
  end
  
endtask
`endif

task read_4_byte;
  regWrEn   = 1'b1;
  #CLKPERIOD;
  #CLKPERIOD;
  #CLKPERIOD;
  #CLKPERIOD;
  regWrEn   = 1'b0;
  regAddr   = 6'h1E;
  #CLKPERIOD;
  $display("%x",regRdData); 
  regAddr   = 6'h1D;
  #CLKPERIOD;
  $display("%x",regRdData); 
  regAddr   = 6'h1C;
  #CLKPERIOD;
  $display("%x",regRdData); 
  regAddr   = 6'h1B;
  #CLKPERIOD;
  $display("%x",regRdData); 
  #CLKPERIOD;
  #CLKPERIOD;
  #CLKPERIOD;
endtask

`ifdef SCAN_EN
task scan_lookup;
integer flop_file;
begin 
   flop_file = $fopen("scan_lu_in.dat","w");
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_33__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_32__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_31__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_30__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_29__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_28__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_27__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_26__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_25__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_24__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_23__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_22__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_21__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_20__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_19__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_18__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_17__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_16__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_15__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_14__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_13__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_12__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_11__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_10__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_9__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_8__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_7__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_6__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_5__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_4__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_3__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_2__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_1__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__319_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__318_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__317_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__316_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__315_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__314_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__313_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__312_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__311_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__310_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__309_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__308_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__307_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__306_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__305_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__304_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__303_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__302_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__301_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__300_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__299_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__298_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__297_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__296_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__295_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__294_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__293_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__292_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__291_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__290_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__289_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__288_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__287_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__286_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__285_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__284_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__283_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__282_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__281_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__280_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__279_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__278_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__277_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__276_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__275_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__274_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__273_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__272_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__271_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__270_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__269_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__268_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__267_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__266_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__265_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__264_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__263_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__262_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__261_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__260_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__259_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__258_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__257_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__256_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__255_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__254_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__253_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__252_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__251_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__250_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__249_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__248_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__247_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__246_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__245_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__244_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__243_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__242_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__241_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__240_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__239_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__238_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__237_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__236_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__235_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__234_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__233_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__232_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__231_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__230_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__229_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__228_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__227_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__226_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__225_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__224_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__223_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__222_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__221_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__220_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__219_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__218_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__217_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__216_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__215_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__214_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__213_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__212_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__211_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__210_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__209_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__208_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__207_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__206_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__205_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__204_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__203_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__202_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__201_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__200_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__199_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__198_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__197_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__196_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__195_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__194_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__193_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__192_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__191_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__190_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__189_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__188_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__187_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__186_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__185_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__184_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__183_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__182_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__181_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__180_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__179_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__178_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__177_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__176_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__175_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__174_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__173_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__172_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__171_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__170_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__169_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__168_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__167_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__166_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__165_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__164_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__163_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__162_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__161_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__160_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__159_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__158_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__157_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__156_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__155_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__154_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__153_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__152_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__151_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__150_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__149_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__148_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__147_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__146_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__145_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__144_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__143_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__142_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__141_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__140_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__139_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__138_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__137_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__136_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__135_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__134_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__133_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__132_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__131_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__130_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__129_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__128_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__127_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__126_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__125_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__124_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__123_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__122_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__121_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__120_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__119_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__118_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__117_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__116_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__115_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__114_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__113_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__112_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__111_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__110_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__109_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__108_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__107_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__106_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__105_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__104_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__103_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__102_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__101_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__100_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__99_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__98_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__97_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__96_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__95_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__94_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__93_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__92_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__91_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__90_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__89_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__88_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__87_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__86_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__85_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__84_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__83_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__82_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__81_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__80_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__79_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__78_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__77_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__76_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__75_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__74_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__73_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__72_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__71_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__70_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__69_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__68_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__67_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__66_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__65_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__64_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__63_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__62_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__61_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__60_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__59_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__58_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__57_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__56_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__55_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__54_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__53_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__52_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__51_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__50_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__49_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__48_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__47_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__46_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__45_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__44_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__43_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__42_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__41_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__40_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__39_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__38_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__37_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__36_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__35_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__34_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__33_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__32_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_0__0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.stallFetch_sync2_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.stallFetch_sync1_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.scratchRegister_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.scratchRegister_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.scratchRegister_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.scratchRegister_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.scratchRegister_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.scratchRegister_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.scratchRegister_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.scratchRegister_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.saluLaneActive_sync_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.saluLaneActive_sync_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.saluLaneActive_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.saluLaneActive_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.saluLaneActive_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.saluLaneActive_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.saluLaneActive_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.rfPartitionActive_sync_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.rfPartitionActive_sync_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.rfPartitionActive_sync_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.rfPartitionActive_sync_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.rfPartitionActive_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.rfPartitionActive_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.rfPartitionActive_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.rfPartitionActive_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.reset_sync2_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.reset_sync1_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.resetFetch_sync2_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.resetFetch_sync1_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.regRdData_o_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.regRdData_o_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.regRdData_o_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.regRdData_o_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.regRdData_o_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.regRdData_o_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.regRdData_o_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.regRdData_o_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.reconfigureCore_sync2_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.reconfigureCore_sync1_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.reconfigDone_latch_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.pipeDrained_latch_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegRun_sync_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegRun_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegGlobalClr_sync_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegGlobalClr_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegData_ioClk_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegClr_sync_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegClr_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegAddr_sync_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegAddr_sync_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegAddr_sync_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegAddr_sync_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegAddr_sync_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegAddr_sync_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegAddr_sync_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegAddr_sync_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegAddr_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegAddr_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegAddr_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegAddr_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegAddr_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegAddr_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegAddr_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.perfMonRegAddr_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.lsqPartitionActive_sync_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.lsqPartitionActive_sync_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.lsqPartitionActive_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.lsqPartitionActive_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.issueLaneActive_sync_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.issueLaneActive_sync_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.issueLaneActive_sync_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.issueLaneActive_sync_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.issueLaneActive_sync_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.issueLaneActive_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.issueLaneActive_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.issueLaneActive_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.issueLaneActive_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.issueLaneActive_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.iqPartitionActive_sync_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.iqPartitionActive_sync_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.iqPartitionActive_sync_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.iqPartitionActive_sync_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.iqPartitionActive_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.iqPartitionActive_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.iqPartitionActive_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.iqPartitionActive_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.instCacheBypass_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrEn_sync_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrEn_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrData_sync_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrData_sync_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrData_sync_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrData_sync_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrData_sync_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrData_sync_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrData_sync_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrData_sync_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrData_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrData_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrData_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrData_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrData_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrData_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrData_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrData_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_sync_reg_10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_sync_reg_9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_sync_reg_8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_sync_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_sync_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_sync_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_sync_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_sync_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_sync_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_sync_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_sync_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_reg_10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_reg_9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_reg_8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchWrAddr_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchRdData_ioClk_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchRdData_ioClk_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchRdData_ioClk_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchRdData_ioClk_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchRdData_ioClk_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchRdData_ioClk_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchRdData_ioClk_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchRdData_ioClk_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchModeEn_sync_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.icScratchModeEn_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.ibuffPartitionActive_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.ibuffPartitionActive_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.ibuffPartitionActive_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.ibuffPartitionActive_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.fetchLaneActive_sync_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.fetchLaneActive_sync_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.fetchLaneActive_sync_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.fetchLaneActive_sync_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.fetchLaneActive_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.fetchLaneActive_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.fetchLaneActive_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.fetchLaneActive_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.execLaneActive_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.execLaneActive_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.execLaneActive_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.execLaneActive_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.execLaneActive_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dispatchLaneActive_sync_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dispatchLaneActive_sync_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dispatchLaneActive_sync_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dispatchLaneActive_sync_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dispatchLaneActive_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dispatchLaneActive_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dispatchLaneActive_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dispatchLaneActive_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrEn_sync_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrEn_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrData_sync_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrData_sync_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrData_sync_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrData_sync_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrData_sync_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrData_sync_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrData_sync_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrData_sync_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrData_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrData_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrData_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrData_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrData_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrData_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrData_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFWrData_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFRdData_ioClk_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFRdData_ioClk_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFRdData_ioClk_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFRdData_ioClk_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFRdData_ioClk_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFRdData_ioClk_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFRdData_ioClk_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFRdData_ioClk_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_sync_reg_8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_sync_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_sync_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_sync_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_sync_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_sync_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_sync_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_sync_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_sync_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_reg_8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugPRFAddr_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTRdData_ioClk_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTRdData_ioClk_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTRdData_ioClk_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTRdData_ioClk_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTRdData_ioClk_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTRdData_ioClk_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTRdData_ioClk_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTAddr_sync_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTAddr_sync_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTAddr_sync_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTAddr_sync_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTAddr_sync_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTAddr_sync_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTAddr_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTAddr_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTAddr_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTAddr_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTAddr_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.debugAMTAddr_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrEn_sync_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrEn_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrData_sync_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrData_sync_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrData_sync_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrData_sync_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrData_sync_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrData_sync_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrData_sync_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrData_sync_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrData_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrData_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrData_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrData_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrData_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrData_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrData_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrData_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_sync_reg_10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_sync_reg_9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_sync_reg_8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_sync_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_sync_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_sync_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_sync_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_sync_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_sync_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_sync_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_sync_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_reg_10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_reg_9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_reg_8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchWrAddr_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchRdData_ioClk_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchRdData_ioClk_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchRdData_ioClk_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchRdData_ioClk_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchRdData_ioClk_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchRdData_ioClk_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchRdData_ioClk_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchRdData_ioClk_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchModeEn_sync_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dcScratchModeEn_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.dataCacheBypass_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_31_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_30_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_29_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_28_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_27_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_26_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_25_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_24_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_23_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_22_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_21_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_20_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_19_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_18_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_17_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_16_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_15_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_14_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_13_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_12_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_11_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_10_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_9_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_8_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_7_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_6_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_5_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.currentInstPC_ioClk_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.commitLaneActive_sync_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.commitLaneActive_sync_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.commitLaneActive_sync_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.commitLaneActive_sync_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.commitLaneActive_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.commitLaneActive_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.commitLaneActive_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.commitLaneActive_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.clearDrainedStatus_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.caluLaneActive_reg_4_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.caluLaneActive_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.caluLaneActive_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.caluLaneActive_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.caluLaneActive_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.cacheModeOverride_sync2_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.cacheModeOverride_sync1_reg.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.alPartitionActive_sync_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.alPartitionActive_sync_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.alPartitionActive_sync_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.alPartitionActive_sync_reg_0_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.alPartitionActive_reg_3_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.alPartitionActive_reg_2_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.alPartitionActive_reg_1_.Q);
$fwrite(flop_file, "%b\n", fab_chip.debCon.alPartitionActive_reg_0_.Q);
end
endtask


task scan_lookup_2;
integer flop_file_2;
begin 
   flop_file_2 = $fopen("scan_lu_in_2.dat","w");
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.valid_array_reg_0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_63__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_62__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_61__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_60__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_59__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_58__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_57__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_56__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_55__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_54__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_53__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_52__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_51__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_50__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_49__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_48__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_47__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_46__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_45__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_44__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_43__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_42__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_41__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_40__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_39__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_38__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_37__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_36__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_35__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_34__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_33__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_32__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_31__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_30__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_29__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_28__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_27__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_26__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_25__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_24__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_23__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_22__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_21__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_20__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_19__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_18__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_17__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_16__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_15__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_14__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_13__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_12__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_11__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_10__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_9__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_8__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_7__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_6__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_5__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_4__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_3__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_2__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_1__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.tag_array_reg_0__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_tag_reg_reg_0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_index_reg_reg_5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_index_reg_reg_4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_index_reg_reg_3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_index_reg_reg_2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_index_reg_reg_1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.pc_index_reg_reg_0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Valid_reg.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Tag_reg_0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Index_reg_5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Index_reg_4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Index_reg_3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Index_reg_2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Index_reg_1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.mshr0Index_reg_0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.miss_d2_reg.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.miss_d1_reg.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrIndex_d1_reg_5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrIndex_d1_reg_4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrIndex_d1_reg_3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrIndex_d1_reg_2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrIndex_d1_reg_1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrIndex_d1_reg_0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrEn_d1_reg.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrData_d1_reg_7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrData_d1_reg_6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrData_d1_reg_5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrData_d1_reg_4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrData_d1_reg_3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrData_d1_reg_2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrData_d1_reg_1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrData_d1_reg_0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrByte_d1_reg_4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrByte_d1_reg_3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrByte_d1_reg_2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrByte_d1_reg_1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchWrByte_d1_reg_0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.icScratchModeEn_d1_reg.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillValid_reg.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillTag_reg_0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillIndex_reg_5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillIndex_reg_4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillIndex_reg_3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillIndex_reg_2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillIndex_reg_1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillIndex_reg_0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.fillData_reg_0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_63__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_62__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_61__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_60__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_59__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_58__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_57__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_56__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_55__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_54__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_53__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_52__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_51__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_50__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_49__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_48__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_47__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_46__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_45__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_44__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_43__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_42__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_41__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_40__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_39__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_38__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_37__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_36__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__62_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__61_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__60_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__59_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__58_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__57_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__56_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__55_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__54_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__53_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__52_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__51_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__50_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__49_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__48_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__47_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__46_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__45_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__44_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__43_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__42_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__41_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__40_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__39_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__38_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__37_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__36_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__35_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__34_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__33_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__32_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__31_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__30_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__29_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__28_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__27_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__26_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__25_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__24_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__23_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__22_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__21_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__20_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__19_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__18_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__17_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__16_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__15_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__14_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__13_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__12_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__11_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__10_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__9_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__8_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__7_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__6_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__5_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__4_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__3_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__2_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__1_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_35__0_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__319_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__318_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__317_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__316_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__315_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__314_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__313_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__312_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__311_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__310_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__309_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__308_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__307_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__306_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__305_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__304_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__303_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__302_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__301_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__300_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__299_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__298_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__297_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__296_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__295_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__294_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__293_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__292_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__291_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__290_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__289_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__288_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__287_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__286_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__285_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__284_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__283_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__282_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__281_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__280_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__279_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__278_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__277_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__276_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__275_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__274_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__273_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__272_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__271_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__270_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__269_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__268_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__267_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__266_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__265_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__264_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__263_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__262_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__261_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__260_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__259_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__258_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__257_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__256_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__255_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__254_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__253_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__252_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__251_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__250_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__249_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__248_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__247_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__246_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__245_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__244_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__243_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__242_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__241_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__240_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__239_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__238_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__237_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__236_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__235_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__234_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__233_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__232_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__231_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__230_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__229_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__228_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__227_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__226_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__225_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__224_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__223_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__222_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__221_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__220_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__219_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__218_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__217_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__216_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__215_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__214_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__213_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__212_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__211_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__210_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__209_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__208_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__207_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__206_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__205_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__204_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__203_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__202_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__201_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__200_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__199_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__198_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__197_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__196_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__195_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__194_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__193_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__192_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__191_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__190_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__189_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__188_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__187_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__186_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__185_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__184_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__183_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__182_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__181_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__180_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__179_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__178_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__177_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__176_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__175_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__174_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__173_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__172_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__171_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__170_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__169_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__168_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__167_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__166_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__165_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__164_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__163_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__162_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__161_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__160_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__159_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__158_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__157_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__156_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__155_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__154_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__153_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__152_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__151_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__150_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__149_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__148_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__147_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__146_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__145_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__144_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__143_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__142_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__141_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__140_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__139_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__138_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__137_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__136_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__135_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__134_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__133_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__132_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__131_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__130_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__129_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__128_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__127_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__126_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__125_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__124_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__123_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__122_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__121_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__120_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__119_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__118_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__117_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__116_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__115_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__114_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__113_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__112_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__111_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__110_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__109_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__108_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__107_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__106_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__105_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__104_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__103_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__102_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__101_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__100_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__99_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__98_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__97_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__96_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__95_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__94_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__93_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__92_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__91_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__90_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__89_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__88_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__87_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__86_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__85_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__84_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__83_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__82_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__81_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__80_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__79_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__78_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__77_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__76_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__75_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__74_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__73_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__72_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__71_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__70_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__69_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__68_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__67_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__66_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__65_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__64_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__63_.Q);
$fwrite(flop_file_2, "%b\n", fab_chip.fabScalar.fs1.l1icache.icache.data_array_reg_34__62_.Q);
end
endtask
`endif
//initial
//begin
////beginConsolidation_reg = 1'b0;
////#(2000*CLKPERIOD);
////stallFetch = 1'b1;
////#(10*CLKPERIOD);
////beginConsolidation_reg = 1'b1;
////#CLKPERIOD;
////beginConsolidation_reg = 1'b0;
//////#(100*CLKPERIOD);
//wait (fabScalar.consolidationDone);
//read_ARF();
//end

//assign fabScalar.beginConsolidation = beginConsolidation_reg;

endmodule
module ANTENNATF(
  input A
  );
endmodule
